
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h96990d7f;
    ram_cell[       1] = 32'h0;  // 32'h74a2cf78;
    ram_cell[       2] = 32'h0;  // 32'h565bffe0;
    ram_cell[       3] = 32'h0;  // 32'h963ceb06;
    ram_cell[       4] = 32'h0;  // 32'hd7db37f6;
    ram_cell[       5] = 32'h0;  // 32'h5aa384af;
    ram_cell[       6] = 32'h0;  // 32'h109b3288;
    ram_cell[       7] = 32'h0;  // 32'h532bd839;
    ram_cell[       8] = 32'h0;  // 32'hac936e5d;
    ram_cell[       9] = 32'h0;  // 32'hc0b498fa;
    ram_cell[      10] = 32'h0;  // 32'h513a1ace;
    ram_cell[      11] = 32'h0;  // 32'h3b060a67;
    ram_cell[      12] = 32'h0;  // 32'h996c7464;
    ram_cell[      13] = 32'h0;  // 32'hd1626e39;
    ram_cell[      14] = 32'h0;  // 32'h0fcf28a7;
    ram_cell[      15] = 32'h0;  // 32'h12bfd9b9;
    ram_cell[      16] = 32'h0;  // 32'h01f3fba7;
    ram_cell[      17] = 32'h0;  // 32'h04757972;
    ram_cell[      18] = 32'h0;  // 32'hf58bf4dd;
    ram_cell[      19] = 32'h0;  // 32'h5c22c924;
    ram_cell[      20] = 32'h0;  // 32'h6a411083;
    ram_cell[      21] = 32'h0;  // 32'h237074a2;
    ram_cell[      22] = 32'h0;  // 32'h4f0d0cc1;
    ram_cell[      23] = 32'h0;  // 32'h6035dac5;
    ram_cell[      24] = 32'h0;  // 32'hc19bb8a2;
    ram_cell[      25] = 32'h0;  // 32'he0321360;
    ram_cell[      26] = 32'h0;  // 32'h1eff4b7c;
    ram_cell[      27] = 32'h0;  // 32'h1c1b78d9;
    ram_cell[      28] = 32'h0;  // 32'hfd9db9cb;
    ram_cell[      29] = 32'h0;  // 32'h9bfdf71d;
    ram_cell[      30] = 32'h0;  // 32'ha7730a7a;
    ram_cell[      31] = 32'h0;  // 32'ha512a4ba;
    ram_cell[      32] = 32'h0;  // 32'hadddd1ec;
    ram_cell[      33] = 32'h0;  // 32'h4e3df057;
    ram_cell[      34] = 32'h0;  // 32'ha3eba29f;
    ram_cell[      35] = 32'h0;  // 32'h84be5ff8;
    ram_cell[      36] = 32'h0;  // 32'ha53a80b8;
    ram_cell[      37] = 32'h0;  // 32'h7e889734;
    ram_cell[      38] = 32'h0;  // 32'hbff3725b;
    ram_cell[      39] = 32'h0;  // 32'hd72569f3;
    ram_cell[      40] = 32'h0;  // 32'h48d1c223;
    ram_cell[      41] = 32'h0;  // 32'h5e15dd68;
    ram_cell[      42] = 32'h0;  // 32'h7f4fb71f;
    ram_cell[      43] = 32'h0;  // 32'hbe7f584a;
    ram_cell[      44] = 32'h0;  // 32'ha14d3c0e;
    ram_cell[      45] = 32'h0;  // 32'h8bb24288;
    ram_cell[      46] = 32'h0;  // 32'h520093a9;
    ram_cell[      47] = 32'h0;  // 32'h901ff38a;
    ram_cell[      48] = 32'h0;  // 32'hcaa36c61;
    ram_cell[      49] = 32'h0;  // 32'hca961c34;
    ram_cell[      50] = 32'h0;  // 32'hf4a43dab;
    ram_cell[      51] = 32'h0;  // 32'h7f96ad2a;
    ram_cell[      52] = 32'h0;  // 32'h595be61a;
    ram_cell[      53] = 32'h0;  // 32'h484ed24a;
    ram_cell[      54] = 32'h0;  // 32'hc72be0d4;
    ram_cell[      55] = 32'h0;  // 32'h801c56e4;
    ram_cell[      56] = 32'h0;  // 32'hb8c6736e;
    ram_cell[      57] = 32'h0;  // 32'h73099e4b;
    ram_cell[      58] = 32'h0;  // 32'hb600d6ee;
    ram_cell[      59] = 32'h0;  // 32'h2358d541;
    ram_cell[      60] = 32'h0;  // 32'h8bccf2ed;
    ram_cell[      61] = 32'h0;  // 32'h675c6b2c;
    ram_cell[      62] = 32'h0;  // 32'ha565d3ae;
    ram_cell[      63] = 32'h0;  // 32'h3c773c98;
    ram_cell[      64] = 32'h0;  // 32'hc6be84e8;
    ram_cell[      65] = 32'h0;  // 32'h805270cf;
    ram_cell[      66] = 32'h0;  // 32'hba167118;
    ram_cell[      67] = 32'h0;  // 32'hf023e588;
    ram_cell[      68] = 32'h0;  // 32'h14e250f5;
    ram_cell[      69] = 32'h0;  // 32'h02a68b4b;
    ram_cell[      70] = 32'h0;  // 32'h68d853b8;
    ram_cell[      71] = 32'h0;  // 32'hc1678d6d;
    ram_cell[      72] = 32'h0;  // 32'h234977f9;
    ram_cell[      73] = 32'h0;  // 32'h22f2b332;
    ram_cell[      74] = 32'h0;  // 32'hd8f272e9;
    ram_cell[      75] = 32'h0;  // 32'h72a7b96a;
    ram_cell[      76] = 32'h0;  // 32'h5a4ff317;
    ram_cell[      77] = 32'h0;  // 32'h0a5c13fd;
    ram_cell[      78] = 32'h0;  // 32'h7a1716d4;
    ram_cell[      79] = 32'h0;  // 32'h88c0964d;
    ram_cell[      80] = 32'h0;  // 32'hbe085f4c;
    ram_cell[      81] = 32'h0;  // 32'hba6868cb;
    ram_cell[      82] = 32'h0;  // 32'h640cb9ad;
    ram_cell[      83] = 32'h0;  // 32'h9e1201e0;
    ram_cell[      84] = 32'h0;  // 32'had473fee;
    ram_cell[      85] = 32'h0;  // 32'h4e584732;
    ram_cell[      86] = 32'h0;  // 32'h4cb44ed6;
    ram_cell[      87] = 32'h0;  // 32'h994740f9;
    ram_cell[      88] = 32'h0;  // 32'h395083a5;
    ram_cell[      89] = 32'h0;  // 32'h225a7dac;
    ram_cell[      90] = 32'h0;  // 32'hf6b40480;
    ram_cell[      91] = 32'h0;  // 32'hcbceee35;
    ram_cell[      92] = 32'h0;  // 32'h4c43bc68;
    ram_cell[      93] = 32'h0;  // 32'h5a9793f4;
    ram_cell[      94] = 32'h0;  // 32'h4405fbd7;
    ram_cell[      95] = 32'h0;  // 32'hecccf879;
    ram_cell[      96] = 32'h0;  // 32'h9d383482;
    ram_cell[      97] = 32'h0;  // 32'hbcc1190b;
    ram_cell[      98] = 32'h0;  // 32'h75935a00;
    ram_cell[      99] = 32'h0;  // 32'hbc1c0a56;
    ram_cell[     100] = 32'h0;  // 32'h3f14f628;
    ram_cell[     101] = 32'h0;  // 32'h0e3ca217;
    ram_cell[     102] = 32'h0;  // 32'h454fed92;
    ram_cell[     103] = 32'h0;  // 32'hda5a01f6;
    ram_cell[     104] = 32'h0;  // 32'h1dab23ef;
    ram_cell[     105] = 32'h0;  // 32'h1b948262;
    ram_cell[     106] = 32'h0;  // 32'h35d3c0e7;
    ram_cell[     107] = 32'h0;  // 32'h97a15a3d;
    ram_cell[     108] = 32'h0;  // 32'h72698858;
    ram_cell[     109] = 32'h0;  // 32'h24d7723b;
    ram_cell[     110] = 32'h0;  // 32'hb8085663;
    ram_cell[     111] = 32'h0;  // 32'h9e9c338f;
    ram_cell[     112] = 32'h0;  // 32'hfa045f1d;
    ram_cell[     113] = 32'h0;  // 32'hb556c218;
    ram_cell[     114] = 32'h0;  // 32'h05ea562a;
    ram_cell[     115] = 32'h0;  // 32'h78f8dcee;
    ram_cell[     116] = 32'h0;  // 32'h2fa7448d;
    ram_cell[     117] = 32'h0;  // 32'h68ab27b2;
    ram_cell[     118] = 32'h0;  // 32'h06ba162b;
    ram_cell[     119] = 32'h0;  // 32'h53453133;
    ram_cell[     120] = 32'h0;  // 32'h4428cb10;
    ram_cell[     121] = 32'h0;  // 32'hc7d69407;
    ram_cell[     122] = 32'h0;  // 32'hd507a077;
    ram_cell[     123] = 32'h0;  // 32'h31efea12;
    ram_cell[     124] = 32'h0;  // 32'h4c6e9870;
    ram_cell[     125] = 32'h0;  // 32'h35724390;
    ram_cell[     126] = 32'h0;  // 32'h857f1af2;
    ram_cell[     127] = 32'h0;  // 32'he8deeb5e;
    ram_cell[     128] = 32'h0;  // 32'h09a93958;
    ram_cell[     129] = 32'h0;  // 32'hc7805bba;
    ram_cell[     130] = 32'h0;  // 32'h4156ecee;
    ram_cell[     131] = 32'h0;  // 32'h82875256;
    ram_cell[     132] = 32'h0;  // 32'hbdb49946;
    ram_cell[     133] = 32'h0;  // 32'hc1f5436f;
    ram_cell[     134] = 32'h0;  // 32'h4ad4338d;
    ram_cell[     135] = 32'h0;  // 32'h4b421e21;
    ram_cell[     136] = 32'h0;  // 32'hbf6249d0;
    ram_cell[     137] = 32'h0;  // 32'hbfba3765;
    ram_cell[     138] = 32'h0;  // 32'hd868695c;
    ram_cell[     139] = 32'h0;  // 32'h968af1d4;
    ram_cell[     140] = 32'h0;  // 32'h6888279f;
    ram_cell[     141] = 32'h0;  // 32'hb87a2d71;
    ram_cell[     142] = 32'h0;  // 32'h57ea2e4f;
    ram_cell[     143] = 32'h0;  // 32'h9f69a5f1;
    ram_cell[     144] = 32'h0;  // 32'h7f96d76e;
    ram_cell[     145] = 32'h0;  // 32'h611e0cdc;
    ram_cell[     146] = 32'h0;  // 32'hd4016996;
    ram_cell[     147] = 32'h0;  // 32'hdca94544;
    ram_cell[     148] = 32'h0;  // 32'hf233ed9b;
    ram_cell[     149] = 32'h0;  // 32'h33e86906;
    ram_cell[     150] = 32'h0;  // 32'ha9d98da1;
    ram_cell[     151] = 32'h0;  // 32'h225b008c;
    ram_cell[     152] = 32'h0;  // 32'h8b79720b;
    ram_cell[     153] = 32'h0;  // 32'h015cde36;
    ram_cell[     154] = 32'h0;  // 32'h2dafc2ff;
    ram_cell[     155] = 32'h0;  // 32'h9efe0217;
    ram_cell[     156] = 32'h0;  // 32'h6bbee798;
    ram_cell[     157] = 32'h0;  // 32'he9c465c3;
    ram_cell[     158] = 32'h0;  // 32'h0da76c30;
    ram_cell[     159] = 32'h0;  // 32'hdd007899;
    ram_cell[     160] = 32'h0;  // 32'h0fe4ab3a;
    ram_cell[     161] = 32'h0;  // 32'h11f17621;
    ram_cell[     162] = 32'h0;  // 32'h9e7dba56;
    ram_cell[     163] = 32'h0;  // 32'h1d1e454d;
    ram_cell[     164] = 32'h0;  // 32'h99248928;
    ram_cell[     165] = 32'h0;  // 32'hf447af42;
    ram_cell[     166] = 32'h0;  // 32'h8aecdf9b;
    ram_cell[     167] = 32'h0;  // 32'h577db764;
    ram_cell[     168] = 32'h0;  // 32'h57b8dca2;
    ram_cell[     169] = 32'h0;  // 32'h07e42acd;
    ram_cell[     170] = 32'h0;  // 32'ha2a698ff;
    ram_cell[     171] = 32'h0;  // 32'hf3746814;
    ram_cell[     172] = 32'h0;  // 32'h2c2ea4e2;
    ram_cell[     173] = 32'h0;  // 32'h18958d33;
    ram_cell[     174] = 32'h0;  // 32'h01088c17;
    ram_cell[     175] = 32'h0;  // 32'h0c58f167;
    ram_cell[     176] = 32'h0;  // 32'h9b9a62d1;
    ram_cell[     177] = 32'h0;  // 32'h5cde780a;
    ram_cell[     178] = 32'h0;  // 32'ha7a9b3bb;
    ram_cell[     179] = 32'h0;  // 32'h300e89f8;
    ram_cell[     180] = 32'h0;  // 32'he6ed0623;
    ram_cell[     181] = 32'h0;  // 32'h3bf21376;
    ram_cell[     182] = 32'h0;  // 32'h530cf92d;
    ram_cell[     183] = 32'h0;  // 32'h14b63bcf;
    ram_cell[     184] = 32'h0;  // 32'h7fd6c51b;
    ram_cell[     185] = 32'h0;  // 32'h7b485a2a;
    ram_cell[     186] = 32'h0;  // 32'h2140c528;
    ram_cell[     187] = 32'h0;  // 32'h1a38037a;
    ram_cell[     188] = 32'h0;  // 32'hda62bbbe;
    ram_cell[     189] = 32'h0;  // 32'h33ca8eb0;
    ram_cell[     190] = 32'h0;  // 32'ha134f2fb;
    ram_cell[     191] = 32'h0;  // 32'h684ecf3e;
    ram_cell[     192] = 32'h0;  // 32'ha634e962;
    ram_cell[     193] = 32'h0;  // 32'ha55466f9;
    ram_cell[     194] = 32'h0;  // 32'h67889213;
    ram_cell[     195] = 32'h0;  // 32'h3695065b;
    ram_cell[     196] = 32'h0;  // 32'h784c8fc4;
    ram_cell[     197] = 32'h0;  // 32'h32d76d91;
    ram_cell[     198] = 32'h0;  // 32'h708f05f0;
    ram_cell[     199] = 32'h0;  // 32'ha80c3dc6;
    ram_cell[     200] = 32'h0;  // 32'ha049dc60;
    ram_cell[     201] = 32'h0;  // 32'hed4a7afd;
    ram_cell[     202] = 32'h0;  // 32'h4afdf3c4;
    ram_cell[     203] = 32'h0;  // 32'h9b4fa8e5;
    ram_cell[     204] = 32'h0;  // 32'h9caeb5f4;
    ram_cell[     205] = 32'h0;  // 32'h7398b97b;
    ram_cell[     206] = 32'h0;  // 32'h8dcce5d2;
    ram_cell[     207] = 32'h0;  // 32'h42cf8148;
    ram_cell[     208] = 32'h0;  // 32'h4ca622ad;
    ram_cell[     209] = 32'h0;  // 32'hb2d12588;
    ram_cell[     210] = 32'h0;  // 32'h496693a6;
    ram_cell[     211] = 32'h0;  // 32'hb6e5e261;
    ram_cell[     212] = 32'h0;  // 32'h53736b09;
    ram_cell[     213] = 32'h0;  // 32'h2fb0058f;
    ram_cell[     214] = 32'h0;  // 32'h7f7320e0;
    ram_cell[     215] = 32'h0;  // 32'h1b7bf54a;
    ram_cell[     216] = 32'h0;  // 32'h6a7259e8;
    ram_cell[     217] = 32'h0;  // 32'h7b3ce4b7;
    ram_cell[     218] = 32'h0;  // 32'h68ab1821;
    ram_cell[     219] = 32'h0;  // 32'hfa7a85ab;
    ram_cell[     220] = 32'h0;  // 32'h631bf127;
    ram_cell[     221] = 32'h0;  // 32'h79a7143a;
    ram_cell[     222] = 32'h0;  // 32'h4b8b009b;
    ram_cell[     223] = 32'h0;  // 32'h1091feb5;
    ram_cell[     224] = 32'h0;  // 32'h7d2d80ff;
    ram_cell[     225] = 32'h0;  // 32'h9d68483c;
    ram_cell[     226] = 32'h0;  // 32'h6c51d801;
    ram_cell[     227] = 32'h0;  // 32'h98aa0c6e;
    ram_cell[     228] = 32'h0;  // 32'hbfcb34df;
    ram_cell[     229] = 32'h0;  // 32'hfee9cf02;
    ram_cell[     230] = 32'h0;  // 32'he17cfdd9;
    ram_cell[     231] = 32'h0;  // 32'h5f73b958;
    ram_cell[     232] = 32'h0;  // 32'h5b200376;
    ram_cell[     233] = 32'h0;  // 32'hd6f1c094;
    ram_cell[     234] = 32'h0;  // 32'hf138f75a;
    ram_cell[     235] = 32'h0;  // 32'h0d68bced;
    ram_cell[     236] = 32'h0;  // 32'h02b3916c;
    ram_cell[     237] = 32'h0;  // 32'h21e031a9;
    ram_cell[     238] = 32'h0;  // 32'h8a3896a3;
    ram_cell[     239] = 32'h0;  // 32'hf2dba5f4;
    ram_cell[     240] = 32'h0;  // 32'hf62f0d7e;
    ram_cell[     241] = 32'h0;  // 32'h3925621d;
    ram_cell[     242] = 32'h0;  // 32'h00e3cb0c;
    ram_cell[     243] = 32'h0;  // 32'hdc4a660d;
    ram_cell[     244] = 32'h0;  // 32'h74068ea1;
    ram_cell[     245] = 32'h0;  // 32'h00e5e1f0;
    ram_cell[     246] = 32'h0;  // 32'h0be0de96;
    ram_cell[     247] = 32'h0;  // 32'h5b88f433;
    ram_cell[     248] = 32'h0;  // 32'ha8a85d1b;
    ram_cell[     249] = 32'h0;  // 32'h93c66ab7;
    ram_cell[     250] = 32'h0;  // 32'ha98ec1e4;
    ram_cell[     251] = 32'h0;  // 32'h4416d483;
    ram_cell[     252] = 32'h0;  // 32'hd9502eec;
    ram_cell[     253] = 32'h0;  // 32'hfbc5fe3e;
    ram_cell[     254] = 32'h0;  // 32'h9e9a22d1;
    ram_cell[     255] = 32'h0;  // 32'hb7ff0103;
    ram_cell[     256] = 32'h0;  // 32'hc2d0b523;
    ram_cell[     257] = 32'h0;  // 32'hb7426285;
    ram_cell[     258] = 32'h0;  // 32'h032b69f2;
    ram_cell[     259] = 32'h0;  // 32'hb641b435;
    ram_cell[     260] = 32'h0;  // 32'h36a90672;
    ram_cell[     261] = 32'h0;  // 32'hce9a65fb;
    ram_cell[     262] = 32'h0;  // 32'h5272747a;
    ram_cell[     263] = 32'h0;  // 32'hbf919637;
    ram_cell[     264] = 32'h0;  // 32'h4bfc323d;
    ram_cell[     265] = 32'h0;  // 32'h9f8f106f;
    ram_cell[     266] = 32'h0;  // 32'h510ec116;
    ram_cell[     267] = 32'h0;  // 32'hd50b2e03;
    ram_cell[     268] = 32'h0;  // 32'hea147199;
    ram_cell[     269] = 32'h0;  // 32'h47e3adf8;
    ram_cell[     270] = 32'h0;  // 32'hd26499a9;
    ram_cell[     271] = 32'h0;  // 32'h595ff9fa;
    ram_cell[     272] = 32'h0;  // 32'he95e9aa7;
    ram_cell[     273] = 32'h0;  // 32'h8c570620;
    ram_cell[     274] = 32'h0;  // 32'he212191f;
    ram_cell[     275] = 32'h0;  // 32'h0737c8d8;
    ram_cell[     276] = 32'h0;  // 32'h5d80ea9a;
    ram_cell[     277] = 32'h0;  // 32'hadf8dfc2;
    ram_cell[     278] = 32'h0;  // 32'h7bbfa1fc;
    ram_cell[     279] = 32'h0;  // 32'h5e271c39;
    ram_cell[     280] = 32'h0;  // 32'h993feaca;
    ram_cell[     281] = 32'h0;  // 32'ha52515ef;
    ram_cell[     282] = 32'h0;  // 32'hd00ab245;
    ram_cell[     283] = 32'h0;  // 32'h691e6197;
    ram_cell[     284] = 32'h0;  // 32'h59ea903f;
    ram_cell[     285] = 32'h0;  // 32'h49ea3edc;
    ram_cell[     286] = 32'h0;  // 32'h7d2a3f42;
    ram_cell[     287] = 32'h0;  // 32'hc209af41;
    ram_cell[     288] = 32'h0;  // 32'h132d29ed;
    ram_cell[     289] = 32'h0;  // 32'headc8897;
    ram_cell[     290] = 32'h0;  // 32'h3bb2ca40;
    ram_cell[     291] = 32'h0;  // 32'hb1fbb310;
    ram_cell[     292] = 32'h0;  // 32'hc69ee571;
    ram_cell[     293] = 32'h0;  // 32'h079bfdde;
    ram_cell[     294] = 32'h0;  // 32'h38cee071;
    ram_cell[     295] = 32'h0;  // 32'h62f5c9dc;
    ram_cell[     296] = 32'h0;  // 32'h866e3c8a;
    ram_cell[     297] = 32'h0;  // 32'h13c871b7;
    ram_cell[     298] = 32'h0;  // 32'ha162c7cb;
    ram_cell[     299] = 32'h0;  // 32'h0053c415;
    ram_cell[     300] = 32'h0;  // 32'ha1b48e59;
    ram_cell[     301] = 32'h0;  // 32'h0411edd3;
    ram_cell[     302] = 32'h0;  // 32'hd45cda0f;
    ram_cell[     303] = 32'h0;  // 32'h3877c5b5;
    ram_cell[     304] = 32'h0;  // 32'hd7b36422;
    ram_cell[     305] = 32'h0;  // 32'h89627aa5;
    ram_cell[     306] = 32'h0;  // 32'h5e092901;
    ram_cell[     307] = 32'h0;  // 32'h6bb30101;
    ram_cell[     308] = 32'h0;  // 32'h4747a479;
    ram_cell[     309] = 32'h0;  // 32'hed73b28a;
    ram_cell[     310] = 32'h0;  // 32'h32ce1fac;
    ram_cell[     311] = 32'h0;  // 32'h31e92532;
    ram_cell[     312] = 32'h0;  // 32'ha5fa1678;
    ram_cell[     313] = 32'h0;  // 32'h9c49566b;
    ram_cell[     314] = 32'h0;  // 32'h64d89adf;
    ram_cell[     315] = 32'h0;  // 32'haa4290ff;
    ram_cell[     316] = 32'h0;  // 32'hcb1cbbd9;
    ram_cell[     317] = 32'h0;  // 32'hdee57847;
    ram_cell[     318] = 32'h0;  // 32'h03f86aa3;
    ram_cell[     319] = 32'h0;  // 32'heaf0818e;
    ram_cell[     320] = 32'h0;  // 32'h33a73556;
    ram_cell[     321] = 32'h0;  // 32'h5ac23f2a;
    ram_cell[     322] = 32'h0;  // 32'h5a9073f8;
    ram_cell[     323] = 32'h0;  // 32'hc9c2760a;
    ram_cell[     324] = 32'h0;  // 32'h7063867d;
    ram_cell[     325] = 32'h0;  // 32'h215c1f21;
    ram_cell[     326] = 32'h0;  // 32'ha8c601bf;
    ram_cell[     327] = 32'h0;  // 32'hf5f16d74;
    ram_cell[     328] = 32'h0;  // 32'hc6228351;
    ram_cell[     329] = 32'h0;  // 32'h823c6d9b;
    ram_cell[     330] = 32'h0;  // 32'h3f9906f9;
    ram_cell[     331] = 32'h0;  // 32'h204a12f7;
    ram_cell[     332] = 32'h0;  // 32'hc51729a6;
    ram_cell[     333] = 32'h0;  // 32'h20ed2281;
    ram_cell[     334] = 32'h0;  // 32'hc0215078;
    ram_cell[     335] = 32'h0;  // 32'hb3dead9f;
    ram_cell[     336] = 32'h0;  // 32'h7f4554a0;
    ram_cell[     337] = 32'h0;  // 32'h544a0a71;
    ram_cell[     338] = 32'h0;  // 32'h12c6892d;
    ram_cell[     339] = 32'h0;  // 32'h3f8596c4;
    ram_cell[     340] = 32'h0;  // 32'h745f655b;
    ram_cell[     341] = 32'h0;  // 32'h27be83df;
    ram_cell[     342] = 32'h0;  // 32'h84d96883;
    ram_cell[     343] = 32'h0;  // 32'he927fadd;
    ram_cell[     344] = 32'h0;  // 32'h8d9c07f4;
    ram_cell[     345] = 32'h0;  // 32'h73c397cc;
    ram_cell[     346] = 32'h0;  // 32'h9f454b3e;
    ram_cell[     347] = 32'h0;  // 32'h00f9618c;
    ram_cell[     348] = 32'h0;  // 32'h4e4b4e6f;
    ram_cell[     349] = 32'h0;  // 32'hfafa2932;
    ram_cell[     350] = 32'h0;  // 32'h47192d5f;
    ram_cell[     351] = 32'h0;  // 32'hbc07ea2e;
    ram_cell[     352] = 32'h0;  // 32'h1ce92eb7;
    ram_cell[     353] = 32'h0;  // 32'h22a1115c;
    ram_cell[     354] = 32'h0;  // 32'h495be591;
    ram_cell[     355] = 32'h0;  // 32'h02c5e0a3;
    ram_cell[     356] = 32'h0;  // 32'ha45bfd26;
    ram_cell[     357] = 32'h0;  // 32'hf794abc2;
    ram_cell[     358] = 32'h0;  // 32'hd3bb401f;
    ram_cell[     359] = 32'h0;  // 32'h86a76b50;
    ram_cell[     360] = 32'h0;  // 32'h31d1d4c6;
    ram_cell[     361] = 32'h0;  // 32'he7d3a476;
    ram_cell[     362] = 32'h0;  // 32'h9fe454b6;
    ram_cell[     363] = 32'h0;  // 32'h54efcfc7;
    ram_cell[     364] = 32'h0;  // 32'h6c98711b;
    ram_cell[     365] = 32'h0;  // 32'hdd5593f8;
    ram_cell[     366] = 32'h0;  // 32'h12cf9a5d;
    ram_cell[     367] = 32'h0;  // 32'h57394082;
    ram_cell[     368] = 32'h0;  // 32'hae4c3b51;
    ram_cell[     369] = 32'h0;  // 32'he4200cbf;
    ram_cell[     370] = 32'h0;  // 32'h41e93e17;
    ram_cell[     371] = 32'h0;  // 32'he008a9cd;
    ram_cell[     372] = 32'h0;  // 32'h33cdf8eb;
    ram_cell[     373] = 32'h0;  // 32'h9789ddc4;
    ram_cell[     374] = 32'h0;  // 32'h577f2f6e;
    ram_cell[     375] = 32'h0;  // 32'hbcd82925;
    ram_cell[     376] = 32'h0;  // 32'h3db41db9;
    ram_cell[     377] = 32'h0;  // 32'h9a6e11f1;
    ram_cell[     378] = 32'h0;  // 32'h140c6884;
    ram_cell[     379] = 32'h0;  // 32'hd0208651;
    ram_cell[     380] = 32'h0;  // 32'h76fcff5e;
    ram_cell[     381] = 32'h0;  // 32'h7050e33a;
    ram_cell[     382] = 32'h0;  // 32'hca345641;
    ram_cell[     383] = 32'h0;  // 32'h19cb90fd;
    ram_cell[     384] = 32'h0;  // 32'h10b68726;
    ram_cell[     385] = 32'h0;  // 32'h76563890;
    ram_cell[     386] = 32'h0;  // 32'h2d4ed011;
    ram_cell[     387] = 32'h0;  // 32'h2783f3f2;
    ram_cell[     388] = 32'h0;  // 32'he8e61002;
    ram_cell[     389] = 32'h0;  // 32'h8c908a40;
    ram_cell[     390] = 32'h0;  // 32'hee43af77;
    ram_cell[     391] = 32'h0;  // 32'h12979f8a;
    ram_cell[     392] = 32'h0;  // 32'h2de5c3fd;
    ram_cell[     393] = 32'h0;  // 32'hc18613ec;
    ram_cell[     394] = 32'h0;  // 32'hc8742353;
    ram_cell[     395] = 32'h0;  // 32'h1ddabfac;
    ram_cell[     396] = 32'h0;  // 32'he5745584;
    ram_cell[     397] = 32'h0;  // 32'h1d4bb797;
    ram_cell[     398] = 32'h0;  // 32'h893ad1d3;
    ram_cell[     399] = 32'h0;  // 32'h5074beb0;
    ram_cell[     400] = 32'h0;  // 32'h04d8bfec;
    ram_cell[     401] = 32'h0;  // 32'h2fa505b3;
    ram_cell[     402] = 32'h0;  // 32'h681cfc2e;
    ram_cell[     403] = 32'h0;  // 32'h4ea8165a;
    ram_cell[     404] = 32'h0;  // 32'h921099ef;
    ram_cell[     405] = 32'h0;  // 32'he3a6405e;
    ram_cell[     406] = 32'h0;  // 32'h43d36270;
    ram_cell[     407] = 32'h0;  // 32'hf9bd2e0d;
    ram_cell[     408] = 32'h0;  // 32'hf858fed4;
    ram_cell[     409] = 32'h0;  // 32'he5539702;
    ram_cell[     410] = 32'h0;  // 32'hee891159;
    ram_cell[     411] = 32'h0;  // 32'h91f9b63f;
    ram_cell[     412] = 32'h0;  // 32'h66bea61b;
    ram_cell[     413] = 32'h0;  // 32'h6a0e0334;
    ram_cell[     414] = 32'h0;  // 32'h7847a939;
    ram_cell[     415] = 32'h0;  // 32'h22fb3cc2;
    ram_cell[     416] = 32'h0;  // 32'hb7fb2937;
    ram_cell[     417] = 32'h0;  // 32'hc77f0a8d;
    ram_cell[     418] = 32'h0;  // 32'h398bdfea;
    ram_cell[     419] = 32'h0;  // 32'haa088b6a;
    ram_cell[     420] = 32'h0;  // 32'h6dc287ab;
    ram_cell[     421] = 32'h0;  // 32'h9ee15f96;
    ram_cell[     422] = 32'h0;  // 32'h79fbb0ca;
    ram_cell[     423] = 32'h0;  // 32'h6b207f2e;
    ram_cell[     424] = 32'h0;  // 32'h76a71024;
    ram_cell[     425] = 32'h0;  // 32'h6d6998bd;
    ram_cell[     426] = 32'h0;  // 32'h6ca27bd1;
    ram_cell[     427] = 32'h0;  // 32'h351ac1c4;
    ram_cell[     428] = 32'h0;  // 32'h0324ac85;
    ram_cell[     429] = 32'h0;  // 32'h39e04806;
    ram_cell[     430] = 32'h0;  // 32'h1bdc7fb3;
    ram_cell[     431] = 32'h0;  // 32'h57dc0421;
    ram_cell[     432] = 32'h0;  // 32'h86990ef7;
    ram_cell[     433] = 32'h0;  // 32'h3387cc63;
    ram_cell[     434] = 32'h0;  // 32'h5b9c75db;
    ram_cell[     435] = 32'h0;  // 32'h5c707a2b;
    ram_cell[     436] = 32'h0;  // 32'h99391e46;
    ram_cell[     437] = 32'h0;  // 32'hb5f6c034;
    ram_cell[     438] = 32'h0;  // 32'he9127d06;
    ram_cell[     439] = 32'h0;  // 32'hd45b2a53;
    ram_cell[     440] = 32'h0;  // 32'h6687535b;
    ram_cell[     441] = 32'h0;  // 32'h4757b67b;
    ram_cell[     442] = 32'h0;  // 32'h359843fe;
    ram_cell[     443] = 32'h0;  // 32'had6763db;
    ram_cell[     444] = 32'h0;  // 32'h84886581;
    ram_cell[     445] = 32'h0;  // 32'hf46f10dc;
    ram_cell[     446] = 32'h0;  // 32'h5ed1a959;
    ram_cell[     447] = 32'h0;  // 32'ha66d944f;
    ram_cell[     448] = 32'h0;  // 32'ha758a3d2;
    ram_cell[     449] = 32'h0;  // 32'hcc543c01;
    ram_cell[     450] = 32'h0;  // 32'h527abf99;
    ram_cell[     451] = 32'h0;  // 32'hebbb8882;
    ram_cell[     452] = 32'h0;  // 32'h27629c0e;
    ram_cell[     453] = 32'h0;  // 32'h5cb5ba75;
    ram_cell[     454] = 32'h0;  // 32'ha6a7bff9;
    ram_cell[     455] = 32'h0;  // 32'h2f7bfe64;
    ram_cell[     456] = 32'h0;  // 32'h4824eba2;
    ram_cell[     457] = 32'h0;  // 32'hf18c9f76;
    ram_cell[     458] = 32'h0;  // 32'h5a382b2c;
    ram_cell[     459] = 32'h0;  // 32'hc72c9d15;
    ram_cell[     460] = 32'h0;  // 32'h95cb7f14;
    ram_cell[     461] = 32'h0;  // 32'hed69cd99;
    ram_cell[     462] = 32'h0;  // 32'h1f7043d3;
    ram_cell[     463] = 32'h0;  // 32'h29d74c5f;
    ram_cell[     464] = 32'h0;  // 32'h13c51bff;
    ram_cell[     465] = 32'h0;  // 32'h2be0d577;
    ram_cell[     466] = 32'h0;  // 32'haa583e76;
    ram_cell[     467] = 32'h0;  // 32'ha0cc447e;
    ram_cell[     468] = 32'h0;  // 32'h432557d8;
    ram_cell[     469] = 32'h0;  // 32'h5f7f1022;
    ram_cell[     470] = 32'h0;  // 32'h463b0b3f;
    ram_cell[     471] = 32'h0;  // 32'h2ac84e4f;
    ram_cell[     472] = 32'h0;  // 32'h5fac3eaf;
    ram_cell[     473] = 32'h0;  // 32'h8d8607bd;
    ram_cell[     474] = 32'h0;  // 32'h3f06ab23;
    ram_cell[     475] = 32'h0;  // 32'he8726688;
    ram_cell[     476] = 32'h0;  // 32'hce4da757;
    ram_cell[     477] = 32'h0;  // 32'h7a71035d;
    ram_cell[     478] = 32'h0;  // 32'hd21e726e;
    ram_cell[     479] = 32'h0;  // 32'hb4cd036c;
    ram_cell[     480] = 32'h0;  // 32'h332cfd50;
    ram_cell[     481] = 32'h0;  // 32'h79365648;
    ram_cell[     482] = 32'h0;  // 32'hd24d4a93;
    ram_cell[     483] = 32'h0;  // 32'h6fc63037;
    ram_cell[     484] = 32'h0;  // 32'h9b6b8aa2;
    ram_cell[     485] = 32'h0;  // 32'h83674931;
    ram_cell[     486] = 32'h0;  // 32'hc47316d7;
    ram_cell[     487] = 32'h0;  // 32'h00466436;
    ram_cell[     488] = 32'h0;  // 32'h145b6e25;
    ram_cell[     489] = 32'h0;  // 32'hf23bde35;
    ram_cell[     490] = 32'h0;  // 32'hcae4883a;
    ram_cell[     491] = 32'h0;  // 32'h633b9caf;
    ram_cell[     492] = 32'h0;  // 32'he5dab494;
    ram_cell[     493] = 32'h0;  // 32'h7fb02afe;
    ram_cell[     494] = 32'h0;  // 32'h94443913;
    ram_cell[     495] = 32'h0;  // 32'h97e5e5b5;
    ram_cell[     496] = 32'h0;  // 32'hf7180c87;
    ram_cell[     497] = 32'h0;  // 32'h58a6c286;
    ram_cell[     498] = 32'h0;  // 32'h58c14edd;
    ram_cell[     499] = 32'h0;  // 32'hd39bf667;
    ram_cell[     500] = 32'h0;  // 32'h9f1a2e9e;
    ram_cell[     501] = 32'h0;  // 32'ha47fd133;
    ram_cell[     502] = 32'h0;  // 32'hcd068ecf;
    ram_cell[     503] = 32'h0;  // 32'hc280cb87;
    ram_cell[     504] = 32'h0;  // 32'hcb567eee;
    ram_cell[     505] = 32'h0;  // 32'hc8c53045;
    ram_cell[     506] = 32'h0;  // 32'h76df4fca;
    ram_cell[     507] = 32'h0;  // 32'h5189f2a4;
    ram_cell[     508] = 32'h0;  // 32'h3a9601c3;
    ram_cell[     509] = 32'h0;  // 32'h445c1b14;
    ram_cell[     510] = 32'h0;  // 32'h46196bf5;
    ram_cell[     511] = 32'h0;  // 32'h8c0442e1;
    ram_cell[     512] = 32'h0;  // 32'h91f5ef16;
    ram_cell[     513] = 32'h0;  // 32'h1c232106;
    ram_cell[     514] = 32'h0;  // 32'he980daf8;
    ram_cell[     515] = 32'h0;  // 32'h05f1dfb2;
    ram_cell[     516] = 32'h0;  // 32'h17bd0c93;
    ram_cell[     517] = 32'h0;  // 32'h502aec56;
    ram_cell[     518] = 32'h0;  // 32'he915dd90;
    ram_cell[     519] = 32'h0;  // 32'h2887f257;
    ram_cell[     520] = 32'h0;  // 32'h4317c2f2;
    ram_cell[     521] = 32'h0;  // 32'h0967dd45;
    ram_cell[     522] = 32'h0;  // 32'hdc6dece8;
    ram_cell[     523] = 32'h0;  // 32'h185406c2;
    ram_cell[     524] = 32'h0;  // 32'h6d488cdb;
    ram_cell[     525] = 32'h0;  // 32'heb181b21;
    ram_cell[     526] = 32'h0;  // 32'hca8b4b7b;
    ram_cell[     527] = 32'h0;  // 32'h5eeaf1be;
    ram_cell[     528] = 32'h0;  // 32'he94696b4;
    ram_cell[     529] = 32'h0;  // 32'h759cb2e0;
    ram_cell[     530] = 32'h0;  // 32'h86383df2;
    ram_cell[     531] = 32'h0;  // 32'h7dab8fbf;
    ram_cell[     532] = 32'h0;  // 32'hdce728d9;
    ram_cell[     533] = 32'h0;  // 32'h81078c42;
    ram_cell[     534] = 32'h0;  // 32'h308e25a0;
    ram_cell[     535] = 32'h0;  // 32'h38ad2e02;
    ram_cell[     536] = 32'h0;  // 32'had2b68a5;
    ram_cell[     537] = 32'h0;  // 32'h753c49db;
    ram_cell[     538] = 32'h0;  // 32'h0d9bccae;
    ram_cell[     539] = 32'h0;  // 32'hb48bfed2;
    ram_cell[     540] = 32'h0;  // 32'he7c674ed;
    ram_cell[     541] = 32'h0;  // 32'h97d1143d;
    ram_cell[     542] = 32'h0;  // 32'h9af26a86;
    ram_cell[     543] = 32'h0;  // 32'hc411ff31;
    ram_cell[     544] = 32'h0;  // 32'h6d89a24f;
    ram_cell[     545] = 32'h0;  // 32'h7ddc6a08;
    ram_cell[     546] = 32'h0;  // 32'h4fdf5be6;
    ram_cell[     547] = 32'h0;  // 32'h1cbf64e4;
    ram_cell[     548] = 32'h0;  // 32'h063ef10e;
    ram_cell[     549] = 32'h0;  // 32'he290bb5c;
    ram_cell[     550] = 32'h0;  // 32'he3384425;
    ram_cell[     551] = 32'h0;  // 32'hf2fd69a7;
    ram_cell[     552] = 32'h0;  // 32'h7815fcf1;
    ram_cell[     553] = 32'h0;  // 32'hf5d0c944;
    ram_cell[     554] = 32'h0;  // 32'h10f447c3;
    ram_cell[     555] = 32'h0;  // 32'ha8d5e60f;
    ram_cell[     556] = 32'h0;  // 32'h312a9c93;
    ram_cell[     557] = 32'h0;  // 32'h64c7aab5;
    ram_cell[     558] = 32'h0;  // 32'h8b9cc0f5;
    ram_cell[     559] = 32'h0;  // 32'hca568f46;
    ram_cell[     560] = 32'h0;  // 32'hd0a83bbc;
    ram_cell[     561] = 32'h0;  // 32'h2fe11321;
    ram_cell[     562] = 32'h0;  // 32'hf0c57dae;
    ram_cell[     563] = 32'h0;  // 32'haaf0870a;
    ram_cell[     564] = 32'h0;  // 32'h09052183;
    ram_cell[     565] = 32'h0;  // 32'ha1fcd7da;
    ram_cell[     566] = 32'h0;  // 32'hddb6eec3;
    ram_cell[     567] = 32'h0;  // 32'h8dbb64de;
    ram_cell[     568] = 32'h0;  // 32'he31b72b9;
    ram_cell[     569] = 32'h0;  // 32'hb72838a8;
    ram_cell[     570] = 32'h0;  // 32'hcca369ff;
    ram_cell[     571] = 32'h0;  // 32'h97dbfa1d;
    ram_cell[     572] = 32'h0;  // 32'hecd72358;
    ram_cell[     573] = 32'h0;  // 32'h27b5495f;
    ram_cell[     574] = 32'h0;  // 32'h8eb28f6f;
    ram_cell[     575] = 32'h0;  // 32'hf6c4a4f1;
    ram_cell[     576] = 32'h0;  // 32'h8e1da83b;
    ram_cell[     577] = 32'h0;  // 32'hfa987e32;
    ram_cell[     578] = 32'h0;  // 32'h36d87fde;
    ram_cell[     579] = 32'h0;  // 32'hd781ddb0;
    ram_cell[     580] = 32'h0;  // 32'hf542d314;
    ram_cell[     581] = 32'h0;  // 32'h6bc13f3c;
    ram_cell[     582] = 32'h0;  // 32'h75e4f773;
    ram_cell[     583] = 32'h0;  // 32'h76a549e3;
    ram_cell[     584] = 32'h0;  // 32'he16adb7f;
    ram_cell[     585] = 32'h0;  // 32'h34d0f962;
    ram_cell[     586] = 32'h0;  // 32'h4f28a26e;
    ram_cell[     587] = 32'h0;  // 32'h1e574c45;
    ram_cell[     588] = 32'h0;  // 32'h49cc1bc0;
    ram_cell[     589] = 32'h0;  // 32'hbb829f23;
    ram_cell[     590] = 32'h0;  // 32'hf7c688e8;
    ram_cell[     591] = 32'h0;  // 32'had7f1633;
    ram_cell[     592] = 32'h0;  // 32'h5a002276;
    ram_cell[     593] = 32'h0;  // 32'h31e4534b;
    ram_cell[     594] = 32'h0;  // 32'h6dabf117;
    ram_cell[     595] = 32'h0;  // 32'h70cae607;
    ram_cell[     596] = 32'h0;  // 32'h839301d5;
    ram_cell[     597] = 32'h0;  // 32'h5c156408;
    ram_cell[     598] = 32'h0;  // 32'hb71a9e72;
    ram_cell[     599] = 32'h0;  // 32'hc45a734d;
    ram_cell[     600] = 32'h0;  // 32'h2d43790d;
    ram_cell[     601] = 32'h0;  // 32'h481caf1a;
    ram_cell[     602] = 32'h0;  // 32'h05e94b2d;
    ram_cell[     603] = 32'h0;  // 32'hddf86c49;
    ram_cell[     604] = 32'h0;  // 32'h0525ce8b;
    ram_cell[     605] = 32'h0;  // 32'h0a37ba09;
    ram_cell[     606] = 32'h0;  // 32'had641568;
    ram_cell[     607] = 32'h0;  // 32'hcd6baf1e;
    ram_cell[     608] = 32'h0;  // 32'h7af7455b;
    ram_cell[     609] = 32'h0;  // 32'hd6bc1803;
    ram_cell[     610] = 32'h0;  // 32'ha14e35b3;
    ram_cell[     611] = 32'h0;  // 32'h703512d2;
    ram_cell[     612] = 32'h0;  // 32'h20e7eedc;
    ram_cell[     613] = 32'h0;  // 32'ha6527c10;
    ram_cell[     614] = 32'h0;  // 32'hd6df9095;
    ram_cell[     615] = 32'h0;  // 32'h3aed5b7c;
    ram_cell[     616] = 32'h0;  // 32'hdd3471e9;
    ram_cell[     617] = 32'h0;  // 32'h8203a91d;
    ram_cell[     618] = 32'h0;  // 32'h21ae1021;
    ram_cell[     619] = 32'h0;  // 32'hf0153429;
    ram_cell[     620] = 32'h0;  // 32'h6b671167;
    ram_cell[     621] = 32'h0;  // 32'h628c2040;
    ram_cell[     622] = 32'h0;  // 32'h9e7288b2;
    ram_cell[     623] = 32'h0;  // 32'h8a27068a;
    ram_cell[     624] = 32'h0;  // 32'h6b479969;
    ram_cell[     625] = 32'h0;  // 32'hce4bf64f;
    ram_cell[     626] = 32'h0;  // 32'he21b4583;
    ram_cell[     627] = 32'h0;  // 32'habed0db4;
    ram_cell[     628] = 32'h0;  // 32'ha8786aef;
    ram_cell[     629] = 32'h0;  // 32'h98c52573;
    ram_cell[     630] = 32'h0;  // 32'h87f509ed;
    ram_cell[     631] = 32'h0;  // 32'h0648b9ba;
    ram_cell[     632] = 32'h0;  // 32'h07250da5;
    ram_cell[     633] = 32'h0;  // 32'h85a1cc31;
    ram_cell[     634] = 32'h0;  // 32'h6136a4a1;
    ram_cell[     635] = 32'h0;  // 32'h1d27ed3a;
    ram_cell[     636] = 32'h0;  // 32'hdbab7d8e;
    ram_cell[     637] = 32'h0;  // 32'h08eee516;
    ram_cell[     638] = 32'h0;  // 32'hf2995043;
    ram_cell[     639] = 32'h0;  // 32'h0f4dd788;
    ram_cell[     640] = 32'h0;  // 32'h4c8716bf;
    ram_cell[     641] = 32'h0;  // 32'h2e711571;
    ram_cell[     642] = 32'h0;  // 32'h7d49501e;
    ram_cell[     643] = 32'h0;  // 32'h8d144724;
    ram_cell[     644] = 32'h0;  // 32'h2adf5c51;
    ram_cell[     645] = 32'h0;  // 32'h4bf6240b;
    ram_cell[     646] = 32'h0;  // 32'haed30fa4;
    ram_cell[     647] = 32'h0;  // 32'h2670ab51;
    ram_cell[     648] = 32'h0;  // 32'ha965534f;
    ram_cell[     649] = 32'h0;  // 32'h5e4d71f4;
    ram_cell[     650] = 32'h0;  // 32'h1495d496;
    ram_cell[     651] = 32'h0;  // 32'h8d83b1b7;
    ram_cell[     652] = 32'h0;  // 32'h2c08cead;
    ram_cell[     653] = 32'h0;  // 32'hf2e028fd;
    ram_cell[     654] = 32'h0;  // 32'ha6a3084e;
    ram_cell[     655] = 32'h0;  // 32'h71931455;
    ram_cell[     656] = 32'h0;  // 32'h3429592a;
    ram_cell[     657] = 32'h0;  // 32'hf0e5b17f;
    ram_cell[     658] = 32'h0;  // 32'hbd3e71c7;
    ram_cell[     659] = 32'h0;  // 32'he01c219d;
    ram_cell[     660] = 32'h0;  // 32'h9f83eb47;
    ram_cell[     661] = 32'h0;  // 32'h78d531b2;
    ram_cell[     662] = 32'h0;  // 32'h637003de;
    ram_cell[     663] = 32'h0;  // 32'h89922077;
    ram_cell[     664] = 32'h0;  // 32'h70d21c8f;
    ram_cell[     665] = 32'h0;  // 32'hbc90cc63;
    ram_cell[     666] = 32'h0;  // 32'h2e704ae5;
    ram_cell[     667] = 32'h0;  // 32'h97a15c23;
    ram_cell[     668] = 32'h0;  // 32'h6b1fe972;
    ram_cell[     669] = 32'h0;  // 32'h9365384c;
    ram_cell[     670] = 32'h0;  // 32'h6dc811ba;
    ram_cell[     671] = 32'h0;  // 32'hbf041139;
    ram_cell[     672] = 32'h0;  // 32'hc1da2bca;
    ram_cell[     673] = 32'h0;  // 32'h13d5f7ec;
    ram_cell[     674] = 32'h0;  // 32'h7a928cd0;
    ram_cell[     675] = 32'h0;  // 32'h1ad7ef31;
    ram_cell[     676] = 32'h0;  // 32'h61153084;
    ram_cell[     677] = 32'h0;  // 32'hb65be3ad;
    ram_cell[     678] = 32'h0;  // 32'h4390a9b7;
    ram_cell[     679] = 32'h0;  // 32'h515d11c0;
    ram_cell[     680] = 32'h0;  // 32'h4b8e90cb;
    ram_cell[     681] = 32'h0;  // 32'h5a88411c;
    ram_cell[     682] = 32'h0;  // 32'h014a3373;
    ram_cell[     683] = 32'h0;  // 32'h6d705502;
    ram_cell[     684] = 32'h0;  // 32'h7a75c1ae;
    ram_cell[     685] = 32'h0;  // 32'h1618718d;
    ram_cell[     686] = 32'h0;  // 32'h3993f95e;
    ram_cell[     687] = 32'h0;  // 32'ha03aaff3;
    ram_cell[     688] = 32'h0;  // 32'hd065737d;
    ram_cell[     689] = 32'h0;  // 32'he9c8d11e;
    ram_cell[     690] = 32'h0;  // 32'h61645347;
    ram_cell[     691] = 32'h0;  // 32'h35a543d5;
    ram_cell[     692] = 32'h0;  // 32'h39873f4c;
    ram_cell[     693] = 32'h0;  // 32'hc01932c5;
    ram_cell[     694] = 32'h0;  // 32'h73d4db47;
    ram_cell[     695] = 32'h0;  // 32'h5346ee44;
    ram_cell[     696] = 32'h0;  // 32'hf923da77;
    ram_cell[     697] = 32'h0;  // 32'h7ca84e95;
    ram_cell[     698] = 32'h0;  // 32'hf1f45b17;
    ram_cell[     699] = 32'h0;  // 32'h2231701c;
    ram_cell[     700] = 32'h0;  // 32'h841ad5a3;
    ram_cell[     701] = 32'h0;  // 32'hc7eb5ec7;
    ram_cell[     702] = 32'h0;  // 32'ha359f38b;
    ram_cell[     703] = 32'h0;  // 32'ha92293ca;
    ram_cell[     704] = 32'h0;  // 32'he45cb8e2;
    ram_cell[     705] = 32'h0;  // 32'h9991a4b2;
    ram_cell[     706] = 32'h0;  // 32'h54fc8e97;
    ram_cell[     707] = 32'h0;  // 32'hb1fc7aa0;
    ram_cell[     708] = 32'h0;  // 32'h400f7021;
    ram_cell[     709] = 32'h0;  // 32'h86c6ace4;
    ram_cell[     710] = 32'h0;  // 32'h4382714d;
    ram_cell[     711] = 32'h0;  // 32'h09e88dfd;
    ram_cell[     712] = 32'h0;  // 32'hd338b95b;
    ram_cell[     713] = 32'h0;  // 32'h188fee42;
    ram_cell[     714] = 32'h0;  // 32'h81ace9e4;
    ram_cell[     715] = 32'h0;  // 32'h95db576a;
    ram_cell[     716] = 32'h0;  // 32'h2c966b3c;
    ram_cell[     717] = 32'h0;  // 32'h566c5952;
    ram_cell[     718] = 32'h0;  // 32'h39aa70d9;
    ram_cell[     719] = 32'h0;  // 32'hda095d59;
    ram_cell[     720] = 32'h0;  // 32'hc29edc06;
    ram_cell[     721] = 32'h0;  // 32'h2471415d;
    ram_cell[     722] = 32'h0;  // 32'h79a231e9;
    ram_cell[     723] = 32'h0;  // 32'h773c3778;
    ram_cell[     724] = 32'h0;  // 32'hcbd446ea;
    ram_cell[     725] = 32'h0;  // 32'hd476be7a;
    ram_cell[     726] = 32'h0;  // 32'he2af47fe;
    ram_cell[     727] = 32'h0;  // 32'hae1caa30;
    ram_cell[     728] = 32'h0;  // 32'hcfb263a6;
    ram_cell[     729] = 32'h0;  // 32'h0148b022;
    ram_cell[     730] = 32'h0;  // 32'hfd75f303;
    ram_cell[     731] = 32'h0;  // 32'h7b9ee9f5;
    ram_cell[     732] = 32'h0;  // 32'h4bb9573c;
    ram_cell[     733] = 32'h0;  // 32'h43492204;
    ram_cell[     734] = 32'h0;  // 32'hc8403274;
    ram_cell[     735] = 32'h0;  // 32'he5710c83;
    ram_cell[     736] = 32'h0;  // 32'hc3010d83;
    ram_cell[     737] = 32'h0;  // 32'h68f68eba;
    ram_cell[     738] = 32'h0;  // 32'hb6065e18;
    ram_cell[     739] = 32'h0;  // 32'h3939b6de;
    ram_cell[     740] = 32'h0;  // 32'h9322eb37;
    ram_cell[     741] = 32'h0;  // 32'ha518e359;
    ram_cell[     742] = 32'h0;  // 32'h1557a8cc;
    ram_cell[     743] = 32'h0;  // 32'h5e8edf20;
    ram_cell[     744] = 32'h0;  // 32'h5f797f47;
    ram_cell[     745] = 32'h0;  // 32'hfd05fd63;
    ram_cell[     746] = 32'h0;  // 32'hb58be9ee;
    ram_cell[     747] = 32'h0;  // 32'h8b3ccc31;
    ram_cell[     748] = 32'h0;  // 32'h0e9f5750;
    ram_cell[     749] = 32'h0;  // 32'hd147b8b7;
    ram_cell[     750] = 32'h0;  // 32'h069808ea;
    ram_cell[     751] = 32'h0;  // 32'h261cc111;
    ram_cell[     752] = 32'h0;  // 32'h489656f8;
    ram_cell[     753] = 32'h0;  // 32'hfaa1e79e;
    ram_cell[     754] = 32'h0;  // 32'h83e8e5c6;
    ram_cell[     755] = 32'h0;  // 32'ha62975d4;
    ram_cell[     756] = 32'h0;  // 32'hb4e75677;
    ram_cell[     757] = 32'h0;  // 32'hc05a6b1a;
    ram_cell[     758] = 32'h0;  // 32'h559c0814;
    ram_cell[     759] = 32'h0;  // 32'h6f872ae7;
    ram_cell[     760] = 32'h0;  // 32'ha7a50a2e;
    ram_cell[     761] = 32'h0;  // 32'h294f017c;
    ram_cell[     762] = 32'h0;  // 32'hb893b4ef;
    ram_cell[     763] = 32'h0;  // 32'h3ed9a42a;
    ram_cell[     764] = 32'h0;  // 32'h772d929f;
    ram_cell[     765] = 32'h0;  // 32'h4b5d89a9;
    ram_cell[     766] = 32'h0;  // 32'h3f23cb12;
    ram_cell[     767] = 32'h0;  // 32'hdeb353e1;
    ram_cell[     768] = 32'h0;  // 32'hcce57231;
    ram_cell[     769] = 32'h0;  // 32'hcfd09db9;
    ram_cell[     770] = 32'h0;  // 32'h15d57395;
    ram_cell[     771] = 32'h0;  // 32'h436e326f;
    ram_cell[     772] = 32'h0;  // 32'h68795754;
    ram_cell[     773] = 32'h0;  // 32'h299bfcaf;
    ram_cell[     774] = 32'h0;  // 32'h86d8ba10;
    ram_cell[     775] = 32'h0;  // 32'h80bc6022;
    ram_cell[     776] = 32'h0;  // 32'h9ae97497;
    ram_cell[     777] = 32'h0;  // 32'ha0fbff16;
    ram_cell[     778] = 32'h0;  // 32'h390b916d;
    ram_cell[     779] = 32'h0;  // 32'h529ad25c;
    ram_cell[     780] = 32'h0;  // 32'h7a274690;
    ram_cell[     781] = 32'h0;  // 32'h6a5c4970;
    ram_cell[     782] = 32'h0;  // 32'h4d9f7cf7;
    ram_cell[     783] = 32'h0;  // 32'h0f47732f;
    ram_cell[     784] = 32'h0;  // 32'h7563f073;
    ram_cell[     785] = 32'h0;  // 32'h1f8b8e86;
    ram_cell[     786] = 32'h0;  // 32'ha62192bf;
    ram_cell[     787] = 32'h0;  // 32'h797510d2;
    ram_cell[     788] = 32'h0;  // 32'h0305b4ec;
    ram_cell[     789] = 32'h0;  // 32'h9a15db38;
    ram_cell[     790] = 32'h0;  // 32'h305f1593;
    ram_cell[     791] = 32'h0;  // 32'h5748b876;
    ram_cell[     792] = 32'h0;  // 32'h66a48f57;
    ram_cell[     793] = 32'h0;  // 32'h8aa4d6c5;
    ram_cell[     794] = 32'h0;  // 32'h1e4be6dc;
    ram_cell[     795] = 32'h0;  // 32'hed13f965;
    ram_cell[     796] = 32'h0;  // 32'h85322ed2;
    ram_cell[     797] = 32'h0;  // 32'h74e52ed2;
    ram_cell[     798] = 32'h0;  // 32'ha0d6347f;
    ram_cell[     799] = 32'h0;  // 32'h07fe4603;
    ram_cell[     800] = 32'h0;  // 32'h5c4e4948;
    ram_cell[     801] = 32'h0;  // 32'h29d5013d;
    ram_cell[     802] = 32'h0;  // 32'hf9457744;
    ram_cell[     803] = 32'h0;  // 32'hdd431513;
    ram_cell[     804] = 32'h0;  // 32'h5221f812;
    ram_cell[     805] = 32'h0;  // 32'h2fa10ecc;
    ram_cell[     806] = 32'h0;  // 32'hf291ebe6;
    ram_cell[     807] = 32'h0;  // 32'h063e793b;
    ram_cell[     808] = 32'h0;  // 32'h59499dc0;
    ram_cell[     809] = 32'h0;  // 32'h112005b1;
    ram_cell[     810] = 32'h0;  // 32'h21b1f16b;
    ram_cell[     811] = 32'h0;  // 32'h1f1fe50b;
    ram_cell[     812] = 32'h0;  // 32'h37b4b012;
    ram_cell[     813] = 32'h0;  // 32'h2ac22b8f;
    ram_cell[     814] = 32'h0;  // 32'h163c8a0b;
    ram_cell[     815] = 32'h0;  // 32'h337907d2;
    ram_cell[     816] = 32'h0;  // 32'h491d8cda;
    ram_cell[     817] = 32'h0;  // 32'h83d5b338;
    ram_cell[     818] = 32'h0;  // 32'hfcb16a15;
    ram_cell[     819] = 32'h0;  // 32'h079f96ef;
    ram_cell[     820] = 32'h0;  // 32'h553081b6;
    ram_cell[     821] = 32'h0;  // 32'h3d667c7b;
    ram_cell[     822] = 32'h0;  // 32'h2454e6d6;
    ram_cell[     823] = 32'h0;  // 32'h7251773d;
    ram_cell[     824] = 32'h0;  // 32'hd7d20d4f;
    ram_cell[     825] = 32'h0;  // 32'hf08d585d;
    ram_cell[     826] = 32'h0;  // 32'h46757153;
    ram_cell[     827] = 32'h0;  // 32'h16c45a7d;
    ram_cell[     828] = 32'h0;  // 32'h6bbad0c0;
    ram_cell[     829] = 32'h0;  // 32'h99098a32;
    ram_cell[     830] = 32'h0;  // 32'h1fc9d67f;
    ram_cell[     831] = 32'h0;  // 32'had087ee7;
    ram_cell[     832] = 32'h0;  // 32'ha97032be;
    ram_cell[     833] = 32'h0;  // 32'hbc38123d;
    ram_cell[     834] = 32'h0;  // 32'h9b1699d8;
    ram_cell[     835] = 32'h0;  // 32'h00847338;
    ram_cell[     836] = 32'h0;  // 32'he8244db7;
    ram_cell[     837] = 32'h0;  // 32'h49d38237;
    ram_cell[     838] = 32'h0;  // 32'hee60b4fe;
    ram_cell[     839] = 32'h0;  // 32'hd1377138;
    ram_cell[     840] = 32'h0;  // 32'h669e5456;
    ram_cell[     841] = 32'h0;  // 32'hf8ff480a;
    ram_cell[     842] = 32'h0;  // 32'hbc7c5494;
    ram_cell[     843] = 32'h0;  // 32'hb1a5e48f;
    ram_cell[     844] = 32'h0;  // 32'h1ad0a57b;
    ram_cell[     845] = 32'h0;  // 32'hcd6bd974;
    ram_cell[     846] = 32'h0;  // 32'hfc2e1bbb;
    ram_cell[     847] = 32'h0;  // 32'h6127a009;
    ram_cell[     848] = 32'h0;  // 32'h90feda5e;
    ram_cell[     849] = 32'h0;  // 32'ha7f19914;
    ram_cell[     850] = 32'h0;  // 32'h46b26dba;
    ram_cell[     851] = 32'h0;  // 32'h291d3c58;
    ram_cell[     852] = 32'h0;  // 32'hc7126c1c;
    ram_cell[     853] = 32'h0;  // 32'h47fbb306;
    ram_cell[     854] = 32'h0;  // 32'hd8de0520;
    ram_cell[     855] = 32'h0;  // 32'h8477ed99;
    ram_cell[     856] = 32'h0;  // 32'h5cb8e685;
    ram_cell[     857] = 32'h0;  // 32'h12e2af02;
    ram_cell[     858] = 32'h0;  // 32'h86c3ae91;
    ram_cell[     859] = 32'h0;  // 32'h0fb35d3c;
    ram_cell[     860] = 32'h0;  // 32'hd7afa2df;
    ram_cell[     861] = 32'h0;  // 32'h47d2edab;
    ram_cell[     862] = 32'h0;  // 32'hfb6c14ff;
    ram_cell[     863] = 32'h0;  // 32'h07f9473b;
    ram_cell[     864] = 32'h0;  // 32'h49968a6b;
    ram_cell[     865] = 32'h0;  // 32'hd467633c;
    ram_cell[     866] = 32'h0;  // 32'ha47eb082;
    ram_cell[     867] = 32'h0;  // 32'h544ba67f;
    ram_cell[     868] = 32'h0;  // 32'hb1bf74db;
    ram_cell[     869] = 32'h0;  // 32'hdb3b27c8;
    ram_cell[     870] = 32'h0;  // 32'hc28e464a;
    ram_cell[     871] = 32'h0;  // 32'hcb021745;
    ram_cell[     872] = 32'h0;  // 32'hb88c47fe;
    ram_cell[     873] = 32'h0;  // 32'hc9b75626;
    ram_cell[     874] = 32'h0;  // 32'h06fc927c;
    ram_cell[     875] = 32'h0;  // 32'h5efb9c4b;
    ram_cell[     876] = 32'h0;  // 32'hb604ea31;
    ram_cell[     877] = 32'h0;  // 32'h2d4475cd;
    ram_cell[     878] = 32'h0;  // 32'h2b1d1aa5;
    ram_cell[     879] = 32'h0;  // 32'h005f565a;
    ram_cell[     880] = 32'h0;  // 32'h6f7a38c9;
    ram_cell[     881] = 32'h0;  // 32'heeef1df7;
    ram_cell[     882] = 32'h0;  // 32'hb9cc0e25;
    ram_cell[     883] = 32'h0;  // 32'haff5182b;
    ram_cell[     884] = 32'h0;  // 32'hbb0f7f5f;
    ram_cell[     885] = 32'h0;  // 32'h172da5f1;
    ram_cell[     886] = 32'h0;  // 32'hf1f1d6b5;
    ram_cell[     887] = 32'h0;  // 32'h0e5bbb56;
    ram_cell[     888] = 32'h0;  // 32'hf515e382;
    ram_cell[     889] = 32'h0;  // 32'hd3dbe484;
    ram_cell[     890] = 32'h0;  // 32'h18cfccee;
    ram_cell[     891] = 32'h0;  // 32'hca91701c;
    ram_cell[     892] = 32'h0;  // 32'h2b430568;
    ram_cell[     893] = 32'h0;  // 32'hf844a9d4;
    ram_cell[     894] = 32'h0;  // 32'hb4c66fa9;
    ram_cell[     895] = 32'h0;  // 32'h8de5ba1a;
    ram_cell[     896] = 32'h0;  // 32'heb9544c0;
    ram_cell[     897] = 32'h0;  // 32'hb6e8367b;
    ram_cell[     898] = 32'h0;  // 32'hd3b6cf84;
    ram_cell[     899] = 32'h0;  // 32'h2162dcce;
    ram_cell[     900] = 32'h0;  // 32'ha4b487a4;
    ram_cell[     901] = 32'h0;  // 32'he0f488a5;
    ram_cell[     902] = 32'h0;  // 32'hd10b2997;
    ram_cell[     903] = 32'h0;  // 32'he867caae;
    ram_cell[     904] = 32'h0;  // 32'h9b544826;
    ram_cell[     905] = 32'h0;  // 32'hfc6c5ec8;
    ram_cell[     906] = 32'h0;  // 32'h5335a1d0;
    ram_cell[     907] = 32'h0;  // 32'hfd4549f8;
    ram_cell[     908] = 32'h0;  // 32'ha479eca1;
    ram_cell[     909] = 32'h0;  // 32'h478efae4;
    ram_cell[     910] = 32'h0;  // 32'hc3e075c2;
    ram_cell[     911] = 32'h0;  // 32'hf05d0fe5;
    ram_cell[     912] = 32'h0;  // 32'hd46df61a;
    ram_cell[     913] = 32'h0;  // 32'h480bc513;
    ram_cell[     914] = 32'h0;  // 32'he5886f7d;
    ram_cell[     915] = 32'h0;  // 32'h1c78f31e;
    ram_cell[     916] = 32'h0;  // 32'he11e3599;
    ram_cell[     917] = 32'h0;  // 32'h73ad7f46;
    ram_cell[     918] = 32'h0;  // 32'h7edd2836;
    ram_cell[     919] = 32'h0;  // 32'h2ce4f024;
    ram_cell[     920] = 32'h0;  // 32'h9f91bfca;
    ram_cell[     921] = 32'h0;  // 32'h26988e27;
    ram_cell[     922] = 32'h0;  // 32'h2955a4f0;
    ram_cell[     923] = 32'h0;  // 32'h4132e678;
    ram_cell[     924] = 32'h0;  // 32'h554f65d7;
    ram_cell[     925] = 32'h0;  // 32'h2c79e9e3;
    ram_cell[     926] = 32'h0;  // 32'h2dcbff27;
    ram_cell[     927] = 32'h0;  // 32'h0ce5119b;
    ram_cell[     928] = 32'h0;  // 32'ha4f63bd9;
    ram_cell[     929] = 32'h0;  // 32'h261aab31;
    ram_cell[     930] = 32'h0;  // 32'h74b66d82;
    ram_cell[     931] = 32'h0;  // 32'hf5670f44;
    ram_cell[     932] = 32'h0;  // 32'hc9e2b7ab;
    ram_cell[     933] = 32'h0;  // 32'h44a242b2;
    ram_cell[     934] = 32'h0;  // 32'hf66f70ab;
    ram_cell[     935] = 32'h0;  // 32'h25ff3804;
    ram_cell[     936] = 32'h0;  // 32'h35dcdac7;
    ram_cell[     937] = 32'h0;  // 32'hd988940c;
    ram_cell[     938] = 32'h0;  // 32'hedcf9615;
    ram_cell[     939] = 32'h0;  // 32'hf82792f2;
    ram_cell[     940] = 32'h0;  // 32'h337a4e57;
    ram_cell[     941] = 32'h0;  // 32'h703f7b6f;
    ram_cell[     942] = 32'h0;  // 32'hc6ec2980;
    ram_cell[     943] = 32'h0;  // 32'h7a9d7ad8;
    ram_cell[     944] = 32'h0;  // 32'h84833da7;
    ram_cell[     945] = 32'h0;  // 32'h8b543105;
    ram_cell[     946] = 32'h0;  // 32'hd540a040;
    ram_cell[     947] = 32'h0;  // 32'h896253e6;
    ram_cell[     948] = 32'h0;  // 32'h80047264;
    ram_cell[     949] = 32'h0;  // 32'hdc482669;
    ram_cell[     950] = 32'h0;  // 32'hbc2c3220;
    ram_cell[     951] = 32'h0;  // 32'hb5741b33;
    ram_cell[     952] = 32'h0;  // 32'h3069f85f;
    ram_cell[     953] = 32'h0;  // 32'he50d3af8;
    ram_cell[     954] = 32'h0;  // 32'h634b8c1d;
    ram_cell[     955] = 32'h0;  // 32'h547eb959;
    ram_cell[     956] = 32'h0;  // 32'hc749cf9a;
    ram_cell[     957] = 32'h0;  // 32'hcbe39c14;
    ram_cell[     958] = 32'h0;  // 32'h12e97473;
    ram_cell[     959] = 32'h0;  // 32'ha0ecd1af;
    ram_cell[     960] = 32'h0;  // 32'hef0abe40;
    ram_cell[     961] = 32'h0;  // 32'h2e9e6d16;
    ram_cell[     962] = 32'h0;  // 32'hba9a258b;
    ram_cell[     963] = 32'h0;  // 32'ha7ca1050;
    ram_cell[     964] = 32'h0;  // 32'ha8ffaa1d;
    ram_cell[     965] = 32'h0;  // 32'h64a0f6c3;
    ram_cell[     966] = 32'h0;  // 32'hf70c721a;
    ram_cell[     967] = 32'h0;  // 32'h10c9465b;
    ram_cell[     968] = 32'h0;  // 32'h3f76f0d5;
    ram_cell[     969] = 32'h0;  // 32'h9c67e76b;
    ram_cell[     970] = 32'h0;  // 32'h6172df39;
    ram_cell[     971] = 32'h0;  // 32'hbec01800;
    ram_cell[     972] = 32'h0;  // 32'h1d11ea90;
    ram_cell[     973] = 32'h0;  // 32'hb69f504c;
    ram_cell[     974] = 32'h0;  // 32'h29f98dc5;
    ram_cell[     975] = 32'h0;  // 32'h509a82e5;
    ram_cell[     976] = 32'h0;  // 32'h34c1323a;
    ram_cell[     977] = 32'h0;  // 32'h3ab67118;
    ram_cell[     978] = 32'h0;  // 32'h8a46c99d;
    ram_cell[     979] = 32'h0;  // 32'h7e4c9cca;
    ram_cell[     980] = 32'h0;  // 32'h85d0987f;
    ram_cell[     981] = 32'h0;  // 32'h67751f42;
    ram_cell[     982] = 32'h0;  // 32'h9a226a56;
    ram_cell[     983] = 32'h0;  // 32'h27daca77;
    ram_cell[     984] = 32'h0;  // 32'h503143cc;
    ram_cell[     985] = 32'h0;  // 32'h8641d1bb;
    ram_cell[     986] = 32'h0;  // 32'h83a10014;
    ram_cell[     987] = 32'h0;  // 32'he78bf0d1;
    ram_cell[     988] = 32'h0;  // 32'ha0de324f;
    ram_cell[     989] = 32'h0;  // 32'h189ee85d;
    ram_cell[     990] = 32'h0;  // 32'h14ef4f99;
    ram_cell[     991] = 32'h0;  // 32'h24353efa;
    ram_cell[     992] = 32'h0;  // 32'hbeabb41b;
    ram_cell[     993] = 32'h0;  // 32'h767757b8;
    ram_cell[     994] = 32'h0;  // 32'h3ecd2e39;
    ram_cell[     995] = 32'h0;  // 32'he6da4834;
    ram_cell[     996] = 32'h0;  // 32'hdc378ba2;
    ram_cell[     997] = 32'h0;  // 32'h96f654db;
    ram_cell[     998] = 32'h0;  // 32'he361ef32;
    ram_cell[     999] = 32'h0;  // 32'h6acf393e;
    ram_cell[    1000] = 32'h0;  // 32'h5702b126;
    ram_cell[    1001] = 32'h0;  // 32'ha9cb9ba2;
    ram_cell[    1002] = 32'h0;  // 32'ha063cee4;
    ram_cell[    1003] = 32'h0;  // 32'h187d2b33;
    ram_cell[    1004] = 32'h0;  // 32'h29f997b6;
    ram_cell[    1005] = 32'h0;  // 32'h56cfe6ae;
    ram_cell[    1006] = 32'h0;  // 32'h09793dd3;
    ram_cell[    1007] = 32'h0;  // 32'h33d443fb;
    ram_cell[    1008] = 32'h0;  // 32'h8bfa50bd;
    ram_cell[    1009] = 32'h0;  // 32'h5c7d648e;
    ram_cell[    1010] = 32'h0;  // 32'hfb854a7c;
    ram_cell[    1011] = 32'h0;  // 32'hd0e7c780;
    ram_cell[    1012] = 32'h0;  // 32'hf285d2ed;
    ram_cell[    1013] = 32'h0;  // 32'h7602666d;
    ram_cell[    1014] = 32'h0;  // 32'h3fecab3f;
    ram_cell[    1015] = 32'h0;  // 32'h93b81d57;
    ram_cell[    1016] = 32'h0;  // 32'hfe0a1bf7;
    ram_cell[    1017] = 32'h0;  // 32'hceb7e5a2;
    ram_cell[    1018] = 32'h0;  // 32'hecbfeba2;
    ram_cell[    1019] = 32'h0;  // 32'h0a8e4d91;
    ram_cell[    1020] = 32'h0;  // 32'h6a370ea4;
    ram_cell[    1021] = 32'h0;  // 32'hf9ad517d;
    ram_cell[    1022] = 32'h0;  // 32'h1f91c9aa;
    ram_cell[    1023] = 32'h0;  // 32'hbdb33df0;
    // src matrix A
    ram_cell[    1024] = 32'he6336a29;
    ram_cell[    1025] = 32'h3c3dbab4;
    ram_cell[    1026] = 32'h16a90308;
    ram_cell[    1027] = 32'h005b7e95;
    ram_cell[    1028] = 32'h33b318b7;
    ram_cell[    1029] = 32'h47bcee2b;
    ram_cell[    1030] = 32'h59e80ae8;
    ram_cell[    1031] = 32'h3a28646d;
    ram_cell[    1032] = 32'h2cd3333a;
    ram_cell[    1033] = 32'h5778a966;
    ram_cell[    1034] = 32'h94c18204;
    ram_cell[    1035] = 32'h39007ae6;
    ram_cell[    1036] = 32'hfc63561d;
    ram_cell[    1037] = 32'h450c1ee2;
    ram_cell[    1038] = 32'h0bfb3d35;
    ram_cell[    1039] = 32'hc03cec36;
    ram_cell[    1040] = 32'hf268b6db;
    ram_cell[    1041] = 32'hf61a39f0;
    ram_cell[    1042] = 32'h420f2fe0;
    ram_cell[    1043] = 32'h014f7ad1;
    ram_cell[    1044] = 32'ha22c9491;
    ram_cell[    1045] = 32'haa97e43a;
    ram_cell[    1046] = 32'hbe0cd5a1;
    ram_cell[    1047] = 32'h27825679;
    ram_cell[    1048] = 32'hef992b62;
    ram_cell[    1049] = 32'hbb103548;
    ram_cell[    1050] = 32'h650bca98;
    ram_cell[    1051] = 32'hc01d125d;
    ram_cell[    1052] = 32'h280bb5a6;
    ram_cell[    1053] = 32'hb90345d0;
    ram_cell[    1054] = 32'h0897bbc8;
    ram_cell[    1055] = 32'hc8323e01;
    ram_cell[    1056] = 32'h8c449f69;
    ram_cell[    1057] = 32'h4d999aea;
    ram_cell[    1058] = 32'h8f49273a;
    ram_cell[    1059] = 32'hda5f662a;
    ram_cell[    1060] = 32'hdd8b30ee;
    ram_cell[    1061] = 32'h9cbf87e3;
    ram_cell[    1062] = 32'hf3846869;
    ram_cell[    1063] = 32'h167ddde3;
    ram_cell[    1064] = 32'hb6c4e5fa;
    ram_cell[    1065] = 32'hb062a4bd;
    ram_cell[    1066] = 32'h03dbbb04;
    ram_cell[    1067] = 32'h8d598dbb;
    ram_cell[    1068] = 32'h73838af8;
    ram_cell[    1069] = 32'h98c169ea;
    ram_cell[    1070] = 32'hdb674da8;
    ram_cell[    1071] = 32'h5b70f859;
    ram_cell[    1072] = 32'hf4760d90;
    ram_cell[    1073] = 32'hab70e1db;
    ram_cell[    1074] = 32'h607a7abc;
    ram_cell[    1075] = 32'he80c6c5c;
    ram_cell[    1076] = 32'h590e64d9;
    ram_cell[    1077] = 32'h30081092;
    ram_cell[    1078] = 32'h777ee18b;
    ram_cell[    1079] = 32'h7c2d9c15;
    ram_cell[    1080] = 32'h8e065b9e;
    ram_cell[    1081] = 32'hc013006c;
    ram_cell[    1082] = 32'h58377cc9;
    ram_cell[    1083] = 32'h1f652507;
    ram_cell[    1084] = 32'h7d848315;
    ram_cell[    1085] = 32'h219bb65b;
    ram_cell[    1086] = 32'h53363940;
    ram_cell[    1087] = 32'hd667b863;
    ram_cell[    1088] = 32'hacd97fdb;
    ram_cell[    1089] = 32'h0da61b05;
    ram_cell[    1090] = 32'ha6c2325f;
    ram_cell[    1091] = 32'h24e4373a;
    ram_cell[    1092] = 32'h77c04312;
    ram_cell[    1093] = 32'hf329e873;
    ram_cell[    1094] = 32'h324bee9f;
    ram_cell[    1095] = 32'h32e748e0;
    ram_cell[    1096] = 32'h52fb0af5;
    ram_cell[    1097] = 32'h3db0faa3;
    ram_cell[    1098] = 32'h98ebc0bc;
    ram_cell[    1099] = 32'h53100d84;
    ram_cell[    1100] = 32'hf50a8548;
    ram_cell[    1101] = 32'heac0611a;
    ram_cell[    1102] = 32'hc2fe4721;
    ram_cell[    1103] = 32'h3c652b77;
    ram_cell[    1104] = 32'h5d6435ac;
    ram_cell[    1105] = 32'h0b7b28fd;
    ram_cell[    1106] = 32'hdbfa9af4;
    ram_cell[    1107] = 32'h4dc91a9f;
    ram_cell[    1108] = 32'h94f641a9;
    ram_cell[    1109] = 32'hf3f3a4e8;
    ram_cell[    1110] = 32'hcb89a309;
    ram_cell[    1111] = 32'h29a871b4;
    ram_cell[    1112] = 32'h030b26a3;
    ram_cell[    1113] = 32'h4c574548;
    ram_cell[    1114] = 32'hd5e4f958;
    ram_cell[    1115] = 32'hdb5121dc;
    ram_cell[    1116] = 32'h5994c134;
    ram_cell[    1117] = 32'h81ed7f4c;
    ram_cell[    1118] = 32'h0dd0fa63;
    ram_cell[    1119] = 32'h2e1e77b9;
    ram_cell[    1120] = 32'h383812be;
    ram_cell[    1121] = 32'hcdf5e474;
    ram_cell[    1122] = 32'h7bad7bf8;
    ram_cell[    1123] = 32'h9db2e3eb;
    ram_cell[    1124] = 32'h5414701f;
    ram_cell[    1125] = 32'h0f0ee28b;
    ram_cell[    1126] = 32'h0c2a80d3;
    ram_cell[    1127] = 32'h85476952;
    ram_cell[    1128] = 32'h415fc61a;
    ram_cell[    1129] = 32'h2d286011;
    ram_cell[    1130] = 32'h469d4158;
    ram_cell[    1131] = 32'h469fe945;
    ram_cell[    1132] = 32'ha6a08c40;
    ram_cell[    1133] = 32'h7e721b48;
    ram_cell[    1134] = 32'h3ea5daa3;
    ram_cell[    1135] = 32'h1abf3746;
    ram_cell[    1136] = 32'h2b1f8bd9;
    ram_cell[    1137] = 32'h7dc9fe56;
    ram_cell[    1138] = 32'h1a76718e;
    ram_cell[    1139] = 32'had9d491b;
    ram_cell[    1140] = 32'ha81e93eb;
    ram_cell[    1141] = 32'hb0359eeb;
    ram_cell[    1142] = 32'h65abbde8;
    ram_cell[    1143] = 32'h8a549ab6;
    ram_cell[    1144] = 32'h781989b5;
    ram_cell[    1145] = 32'h6ab3e343;
    ram_cell[    1146] = 32'h0456356c;
    ram_cell[    1147] = 32'h9f4e58df;
    ram_cell[    1148] = 32'h5812a5d6;
    ram_cell[    1149] = 32'h8ee0c4d1;
    ram_cell[    1150] = 32'h48edf2f7;
    ram_cell[    1151] = 32'h3ca6fc35;
    ram_cell[    1152] = 32'h2ac40361;
    ram_cell[    1153] = 32'h65d3c80f;
    ram_cell[    1154] = 32'h9f3cff6f;
    ram_cell[    1155] = 32'h8d36ef62;
    ram_cell[    1156] = 32'hbc24ee6b;
    ram_cell[    1157] = 32'hb779d5d5;
    ram_cell[    1158] = 32'hf513f86c;
    ram_cell[    1159] = 32'hb2a77c60;
    ram_cell[    1160] = 32'hd3668a53;
    ram_cell[    1161] = 32'hbbbb9788;
    ram_cell[    1162] = 32'h7cf8ca21;
    ram_cell[    1163] = 32'hd4d7183a;
    ram_cell[    1164] = 32'h25360353;
    ram_cell[    1165] = 32'h8e34a3d7;
    ram_cell[    1166] = 32'h5b7a3838;
    ram_cell[    1167] = 32'hfa1f51b4;
    ram_cell[    1168] = 32'h6959559f;
    ram_cell[    1169] = 32'hc8221afd;
    ram_cell[    1170] = 32'hd7810a14;
    ram_cell[    1171] = 32'hdea1a42d;
    ram_cell[    1172] = 32'h577de3b5;
    ram_cell[    1173] = 32'h44452e1f;
    ram_cell[    1174] = 32'h71ab5150;
    ram_cell[    1175] = 32'h98f3651b;
    ram_cell[    1176] = 32'h477d2fef;
    ram_cell[    1177] = 32'hd0f75a25;
    ram_cell[    1178] = 32'h793553a6;
    ram_cell[    1179] = 32'hdb28fd9a;
    ram_cell[    1180] = 32'hcd412518;
    ram_cell[    1181] = 32'hc976d2e1;
    ram_cell[    1182] = 32'he8cfc2e7;
    ram_cell[    1183] = 32'he1616034;
    ram_cell[    1184] = 32'h34232a64;
    ram_cell[    1185] = 32'h055c6a37;
    ram_cell[    1186] = 32'h91fa9125;
    ram_cell[    1187] = 32'hf6593254;
    ram_cell[    1188] = 32'h5574f7f1;
    ram_cell[    1189] = 32'hf2ee4d2f;
    ram_cell[    1190] = 32'h4c29619b;
    ram_cell[    1191] = 32'hde1cdc21;
    ram_cell[    1192] = 32'h13b5fa6e;
    ram_cell[    1193] = 32'hb728783d;
    ram_cell[    1194] = 32'h36354fec;
    ram_cell[    1195] = 32'h28f6f43a;
    ram_cell[    1196] = 32'h5be53a99;
    ram_cell[    1197] = 32'hbb89300d;
    ram_cell[    1198] = 32'h7f920dd6;
    ram_cell[    1199] = 32'hf5df65fe;
    ram_cell[    1200] = 32'hf63afed6;
    ram_cell[    1201] = 32'h5dcdcd5c;
    ram_cell[    1202] = 32'hb0e67fc8;
    ram_cell[    1203] = 32'h67c71049;
    ram_cell[    1204] = 32'hb1df9d91;
    ram_cell[    1205] = 32'hec82fbd4;
    ram_cell[    1206] = 32'h21f7f3ef;
    ram_cell[    1207] = 32'hed1e9577;
    ram_cell[    1208] = 32'hd17354e1;
    ram_cell[    1209] = 32'hd791eaa5;
    ram_cell[    1210] = 32'h81d6a4e5;
    ram_cell[    1211] = 32'hd1d95e48;
    ram_cell[    1212] = 32'h4445a3d4;
    ram_cell[    1213] = 32'h76a2de59;
    ram_cell[    1214] = 32'hd171930d;
    ram_cell[    1215] = 32'hc609706c;
    ram_cell[    1216] = 32'h2c778e58;
    ram_cell[    1217] = 32'h4f2a9615;
    ram_cell[    1218] = 32'h7f66b412;
    ram_cell[    1219] = 32'h5687d1ee;
    ram_cell[    1220] = 32'h46118d2b;
    ram_cell[    1221] = 32'hfe2f4ad8;
    ram_cell[    1222] = 32'hfb646baa;
    ram_cell[    1223] = 32'hf537899c;
    ram_cell[    1224] = 32'h7c100a95;
    ram_cell[    1225] = 32'h385a1479;
    ram_cell[    1226] = 32'h6fc77176;
    ram_cell[    1227] = 32'h052d5650;
    ram_cell[    1228] = 32'h6bcf3355;
    ram_cell[    1229] = 32'h92c82d72;
    ram_cell[    1230] = 32'hbd184e1f;
    ram_cell[    1231] = 32'h6c604ee4;
    ram_cell[    1232] = 32'ha842c437;
    ram_cell[    1233] = 32'h25e47fe2;
    ram_cell[    1234] = 32'h76e54c17;
    ram_cell[    1235] = 32'h6a28baf1;
    ram_cell[    1236] = 32'h0096878d;
    ram_cell[    1237] = 32'h4346e09c;
    ram_cell[    1238] = 32'h1c9d0afd;
    ram_cell[    1239] = 32'hab211b3f;
    ram_cell[    1240] = 32'h68f6e5c8;
    ram_cell[    1241] = 32'he2d20921;
    ram_cell[    1242] = 32'h7563e395;
    ram_cell[    1243] = 32'hd4cf2e5b;
    ram_cell[    1244] = 32'h9fcdd892;
    ram_cell[    1245] = 32'h8bd07503;
    ram_cell[    1246] = 32'h2d1581cf;
    ram_cell[    1247] = 32'h67056c38;
    ram_cell[    1248] = 32'hd90fa8b8;
    ram_cell[    1249] = 32'h1742e24c;
    ram_cell[    1250] = 32'hf2004295;
    ram_cell[    1251] = 32'h174b4e93;
    ram_cell[    1252] = 32'ha8e63c0c;
    ram_cell[    1253] = 32'h323ad1af;
    ram_cell[    1254] = 32'h7e0fcbff;
    ram_cell[    1255] = 32'h595270f9;
    ram_cell[    1256] = 32'h8b9afafd;
    ram_cell[    1257] = 32'hd105b8bf;
    ram_cell[    1258] = 32'hd903c43c;
    ram_cell[    1259] = 32'h67eaf29f;
    ram_cell[    1260] = 32'h3e9c5b23;
    ram_cell[    1261] = 32'h9f11ae8d;
    ram_cell[    1262] = 32'h336c8c45;
    ram_cell[    1263] = 32'h9a810b01;
    ram_cell[    1264] = 32'h6463e562;
    ram_cell[    1265] = 32'h5d420dd5;
    ram_cell[    1266] = 32'h2789a748;
    ram_cell[    1267] = 32'h31622e3b;
    ram_cell[    1268] = 32'hf5613ee2;
    ram_cell[    1269] = 32'hc3d1ff96;
    ram_cell[    1270] = 32'hbc558601;
    ram_cell[    1271] = 32'h608f43c7;
    ram_cell[    1272] = 32'h79024c9b;
    ram_cell[    1273] = 32'h02b18ed3;
    ram_cell[    1274] = 32'h12d0a8dd;
    ram_cell[    1275] = 32'h559add0f;
    ram_cell[    1276] = 32'h46c0bb1b;
    ram_cell[    1277] = 32'hb35f319c;
    ram_cell[    1278] = 32'h0e0be4d6;
    ram_cell[    1279] = 32'h23d9b256;
    ram_cell[    1280] = 32'h94326cf8;
    ram_cell[    1281] = 32'haf8001e5;
    ram_cell[    1282] = 32'h7e19a268;
    ram_cell[    1283] = 32'h4433f61c;
    ram_cell[    1284] = 32'haee361c2;
    ram_cell[    1285] = 32'h0dc47891;
    ram_cell[    1286] = 32'h3ca0914b;
    ram_cell[    1287] = 32'h5d86d365;
    ram_cell[    1288] = 32'hc54f1bf9;
    ram_cell[    1289] = 32'h0d5bb67b;
    ram_cell[    1290] = 32'hd02aab58;
    ram_cell[    1291] = 32'h1b700553;
    ram_cell[    1292] = 32'h76eb0540;
    ram_cell[    1293] = 32'he1b39dc1;
    ram_cell[    1294] = 32'h4926192d;
    ram_cell[    1295] = 32'hffece363;
    ram_cell[    1296] = 32'h8b81424d;
    ram_cell[    1297] = 32'h27335dfa;
    ram_cell[    1298] = 32'h13161eec;
    ram_cell[    1299] = 32'h85c3b626;
    ram_cell[    1300] = 32'h2c8f6296;
    ram_cell[    1301] = 32'h8e45c8df;
    ram_cell[    1302] = 32'hacae241c;
    ram_cell[    1303] = 32'h66a0ea86;
    ram_cell[    1304] = 32'hfecc5e41;
    ram_cell[    1305] = 32'h891a6490;
    ram_cell[    1306] = 32'h31a672b3;
    ram_cell[    1307] = 32'h4918005d;
    ram_cell[    1308] = 32'hb4814603;
    ram_cell[    1309] = 32'haca99715;
    ram_cell[    1310] = 32'hdbc329fa;
    ram_cell[    1311] = 32'h70e1ab6c;
    ram_cell[    1312] = 32'h4bb95fa3;
    ram_cell[    1313] = 32'ha932e9ca;
    ram_cell[    1314] = 32'h6a2ccc8f;
    ram_cell[    1315] = 32'h7de506dc;
    ram_cell[    1316] = 32'hbc965434;
    ram_cell[    1317] = 32'h5cc6df2b;
    ram_cell[    1318] = 32'h56bede2a;
    ram_cell[    1319] = 32'h57273662;
    ram_cell[    1320] = 32'h826c28a8;
    ram_cell[    1321] = 32'h7a35aace;
    ram_cell[    1322] = 32'h284938bc;
    ram_cell[    1323] = 32'h1f3741f0;
    ram_cell[    1324] = 32'h522c61a7;
    ram_cell[    1325] = 32'h95ba7bae;
    ram_cell[    1326] = 32'h051cb55b;
    ram_cell[    1327] = 32'he65a8423;
    ram_cell[    1328] = 32'hd1b610c4;
    ram_cell[    1329] = 32'h7adcfa25;
    ram_cell[    1330] = 32'hf85a0657;
    ram_cell[    1331] = 32'h773d39c6;
    ram_cell[    1332] = 32'h1ef3e721;
    ram_cell[    1333] = 32'h2d0d6ad5;
    ram_cell[    1334] = 32'haf5eff0b;
    ram_cell[    1335] = 32'he9ec9e1d;
    ram_cell[    1336] = 32'hda271f10;
    ram_cell[    1337] = 32'hdb5b7988;
    ram_cell[    1338] = 32'h61c00776;
    ram_cell[    1339] = 32'h1ea34057;
    ram_cell[    1340] = 32'h2b5434a2;
    ram_cell[    1341] = 32'h5c549c80;
    ram_cell[    1342] = 32'hdb60c2b8;
    ram_cell[    1343] = 32'heca54287;
    ram_cell[    1344] = 32'h2268108f;
    ram_cell[    1345] = 32'hcef974d0;
    ram_cell[    1346] = 32'h20dd55fb;
    ram_cell[    1347] = 32'hd2a9bbfd;
    ram_cell[    1348] = 32'hf30e02ba;
    ram_cell[    1349] = 32'h124ac879;
    ram_cell[    1350] = 32'h55b8b334;
    ram_cell[    1351] = 32'h052ec722;
    ram_cell[    1352] = 32'ha66d46f6;
    ram_cell[    1353] = 32'hb6b6f757;
    ram_cell[    1354] = 32'h4b5e7bff;
    ram_cell[    1355] = 32'h079827e1;
    ram_cell[    1356] = 32'h0136e8bc;
    ram_cell[    1357] = 32'h8a7436c7;
    ram_cell[    1358] = 32'h166f9a7d;
    ram_cell[    1359] = 32'hc6d83a50;
    ram_cell[    1360] = 32'he63de1cb;
    ram_cell[    1361] = 32'h4389040a;
    ram_cell[    1362] = 32'ha3d603fd;
    ram_cell[    1363] = 32'h333bc603;
    ram_cell[    1364] = 32'hdd3ef6c2;
    ram_cell[    1365] = 32'hae6dec06;
    ram_cell[    1366] = 32'hf85e0bb1;
    ram_cell[    1367] = 32'h9b2bb638;
    ram_cell[    1368] = 32'h67429a9a;
    ram_cell[    1369] = 32'h4eb5eaac;
    ram_cell[    1370] = 32'h9a396687;
    ram_cell[    1371] = 32'hd34e71db;
    ram_cell[    1372] = 32'hc39cb682;
    ram_cell[    1373] = 32'hcbc21bcc;
    ram_cell[    1374] = 32'h313300b8;
    ram_cell[    1375] = 32'hf1820d66;
    ram_cell[    1376] = 32'he07eabc9;
    ram_cell[    1377] = 32'h0a29c372;
    ram_cell[    1378] = 32'h3cbc55e7;
    ram_cell[    1379] = 32'hb45c2325;
    ram_cell[    1380] = 32'h0b2b33f6;
    ram_cell[    1381] = 32'h038124ec;
    ram_cell[    1382] = 32'h0b8bd3f1;
    ram_cell[    1383] = 32'h5cd3d37d;
    ram_cell[    1384] = 32'hc94326b4;
    ram_cell[    1385] = 32'h7b0a6de6;
    ram_cell[    1386] = 32'h62cd05af;
    ram_cell[    1387] = 32'h82306db2;
    ram_cell[    1388] = 32'h355fd197;
    ram_cell[    1389] = 32'h9248a03d;
    ram_cell[    1390] = 32'h96fe424d;
    ram_cell[    1391] = 32'hc01740de;
    ram_cell[    1392] = 32'hbf0db378;
    ram_cell[    1393] = 32'h4111c694;
    ram_cell[    1394] = 32'h8ce261be;
    ram_cell[    1395] = 32'h780ab111;
    ram_cell[    1396] = 32'h31dca1fb;
    ram_cell[    1397] = 32'hfb138d68;
    ram_cell[    1398] = 32'h2a0c5f94;
    ram_cell[    1399] = 32'hfedb9bc2;
    ram_cell[    1400] = 32'h5f63a3bb;
    ram_cell[    1401] = 32'h50f125d1;
    ram_cell[    1402] = 32'h21290db7;
    ram_cell[    1403] = 32'h87a72aea;
    ram_cell[    1404] = 32'h55a2932d;
    ram_cell[    1405] = 32'h5d505409;
    ram_cell[    1406] = 32'h3ef6a365;
    ram_cell[    1407] = 32'hba8fe7f9;
    ram_cell[    1408] = 32'h71cd02c3;
    ram_cell[    1409] = 32'h0b44d018;
    ram_cell[    1410] = 32'h2df44790;
    ram_cell[    1411] = 32'h4ada8afc;
    ram_cell[    1412] = 32'h49c71789;
    ram_cell[    1413] = 32'hf807c91e;
    ram_cell[    1414] = 32'hb9811134;
    ram_cell[    1415] = 32'h8336629e;
    ram_cell[    1416] = 32'h7d210b25;
    ram_cell[    1417] = 32'h0b07e321;
    ram_cell[    1418] = 32'hdd82e974;
    ram_cell[    1419] = 32'h59358eaf;
    ram_cell[    1420] = 32'h2875ec2d;
    ram_cell[    1421] = 32'h981e154d;
    ram_cell[    1422] = 32'he22c5743;
    ram_cell[    1423] = 32'h3a9a9866;
    ram_cell[    1424] = 32'hb76b11dd;
    ram_cell[    1425] = 32'hb8fe0a65;
    ram_cell[    1426] = 32'h0037b036;
    ram_cell[    1427] = 32'h9cca277b;
    ram_cell[    1428] = 32'h51b3dfd9;
    ram_cell[    1429] = 32'h50b2d454;
    ram_cell[    1430] = 32'hb060f4a1;
    ram_cell[    1431] = 32'hb5bdbb75;
    ram_cell[    1432] = 32'hd1b2ae9b;
    ram_cell[    1433] = 32'h72cac177;
    ram_cell[    1434] = 32'hdca5fc5e;
    ram_cell[    1435] = 32'hc8757911;
    ram_cell[    1436] = 32'h02db5272;
    ram_cell[    1437] = 32'h18a856e7;
    ram_cell[    1438] = 32'h90dfb0cb;
    ram_cell[    1439] = 32'h368e9f83;
    ram_cell[    1440] = 32'hf4ad7205;
    ram_cell[    1441] = 32'h4c85c76d;
    ram_cell[    1442] = 32'h4fd48563;
    ram_cell[    1443] = 32'h2780f3cd;
    ram_cell[    1444] = 32'ha2060161;
    ram_cell[    1445] = 32'h6428c3e5;
    ram_cell[    1446] = 32'h9322031e;
    ram_cell[    1447] = 32'h9d6748a4;
    ram_cell[    1448] = 32'habb65c8a;
    ram_cell[    1449] = 32'h5bcda72e;
    ram_cell[    1450] = 32'h5d2a86e6;
    ram_cell[    1451] = 32'h202ec4a4;
    ram_cell[    1452] = 32'h5bd68df6;
    ram_cell[    1453] = 32'h8b0caacb;
    ram_cell[    1454] = 32'h4966e87c;
    ram_cell[    1455] = 32'heb87e90e;
    ram_cell[    1456] = 32'h90a224a0;
    ram_cell[    1457] = 32'h3889928f;
    ram_cell[    1458] = 32'h3b5b9f2d;
    ram_cell[    1459] = 32'h9a530dbf;
    ram_cell[    1460] = 32'h1e5de611;
    ram_cell[    1461] = 32'h8d3a6f3c;
    ram_cell[    1462] = 32'h4fd3b40c;
    ram_cell[    1463] = 32'hc3f3ce80;
    ram_cell[    1464] = 32'h2e1a35c1;
    ram_cell[    1465] = 32'h8bc2d9b1;
    ram_cell[    1466] = 32'h6cc5a40e;
    ram_cell[    1467] = 32'ha9856708;
    ram_cell[    1468] = 32'h6cf3f101;
    ram_cell[    1469] = 32'hce15dd4e;
    ram_cell[    1470] = 32'hc9b3992d;
    ram_cell[    1471] = 32'ha46dfe63;
    ram_cell[    1472] = 32'hefa8f64d;
    ram_cell[    1473] = 32'h9f97a903;
    ram_cell[    1474] = 32'h255af7a5;
    ram_cell[    1475] = 32'h3d89595e;
    ram_cell[    1476] = 32'h27eee14a;
    ram_cell[    1477] = 32'h295f9d8a;
    ram_cell[    1478] = 32'h3b8c6fc3;
    ram_cell[    1479] = 32'hf75b9382;
    ram_cell[    1480] = 32'h1f77ec61;
    ram_cell[    1481] = 32'hf38fd5c3;
    ram_cell[    1482] = 32'hef1c4873;
    ram_cell[    1483] = 32'hd173682b;
    ram_cell[    1484] = 32'h74e2c1fa;
    ram_cell[    1485] = 32'h46414079;
    ram_cell[    1486] = 32'h4f40965e;
    ram_cell[    1487] = 32'hd7b1bd3e;
    ram_cell[    1488] = 32'heaab60fa;
    ram_cell[    1489] = 32'h9a351aca;
    ram_cell[    1490] = 32'he9db214e;
    ram_cell[    1491] = 32'h10a4fe1b;
    ram_cell[    1492] = 32'hdc6869ae;
    ram_cell[    1493] = 32'hb6ba9df8;
    ram_cell[    1494] = 32'h86597e7a;
    ram_cell[    1495] = 32'hdd999fa8;
    ram_cell[    1496] = 32'h70073620;
    ram_cell[    1497] = 32'hee7f6293;
    ram_cell[    1498] = 32'hf5e2b0e9;
    ram_cell[    1499] = 32'h01bd25f9;
    ram_cell[    1500] = 32'hf5472d60;
    ram_cell[    1501] = 32'hac003724;
    ram_cell[    1502] = 32'h5500e4c4;
    ram_cell[    1503] = 32'hb9c04276;
    ram_cell[    1504] = 32'h6703a2f3;
    ram_cell[    1505] = 32'hf192b8d1;
    ram_cell[    1506] = 32'hf96e9ccb;
    ram_cell[    1507] = 32'h93b0b4b3;
    ram_cell[    1508] = 32'hce1a4221;
    ram_cell[    1509] = 32'h8c7e81cb;
    ram_cell[    1510] = 32'h26fe66ed;
    ram_cell[    1511] = 32'h8cebf895;
    ram_cell[    1512] = 32'hbc75e893;
    ram_cell[    1513] = 32'h5bcfeff2;
    ram_cell[    1514] = 32'h9a4d60ba;
    ram_cell[    1515] = 32'h04218709;
    ram_cell[    1516] = 32'hdc832b9d;
    ram_cell[    1517] = 32'h3ce405c4;
    ram_cell[    1518] = 32'h7c0dc95e;
    ram_cell[    1519] = 32'h4616329a;
    ram_cell[    1520] = 32'h060f3997;
    ram_cell[    1521] = 32'h0684adc6;
    ram_cell[    1522] = 32'hd2e8715d;
    ram_cell[    1523] = 32'he974c94c;
    ram_cell[    1524] = 32'h469e2a3d;
    ram_cell[    1525] = 32'h4db50b40;
    ram_cell[    1526] = 32'h5221ea66;
    ram_cell[    1527] = 32'h12455071;
    ram_cell[    1528] = 32'hf38d263f;
    ram_cell[    1529] = 32'h608705e3;
    ram_cell[    1530] = 32'hd93e0982;
    ram_cell[    1531] = 32'h2e118120;
    ram_cell[    1532] = 32'h9b7fbb60;
    ram_cell[    1533] = 32'he90447f0;
    ram_cell[    1534] = 32'heb6ef934;
    ram_cell[    1535] = 32'h17bada99;
    ram_cell[    1536] = 32'haafec13d;
    ram_cell[    1537] = 32'h6f499b95;
    ram_cell[    1538] = 32'h7e916387;
    ram_cell[    1539] = 32'hbfc3dad6;
    ram_cell[    1540] = 32'hc2508af4;
    ram_cell[    1541] = 32'hd9b7e920;
    ram_cell[    1542] = 32'ha67495a1;
    ram_cell[    1543] = 32'hf53f8dbf;
    ram_cell[    1544] = 32'h99592053;
    ram_cell[    1545] = 32'h94e23b6a;
    ram_cell[    1546] = 32'h007e2e5d;
    ram_cell[    1547] = 32'hee94e611;
    ram_cell[    1548] = 32'hba630f7b;
    ram_cell[    1549] = 32'hf28dad14;
    ram_cell[    1550] = 32'h292083dc;
    ram_cell[    1551] = 32'h85833bdd;
    ram_cell[    1552] = 32'had1f0a2a;
    ram_cell[    1553] = 32'ha829be11;
    ram_cell[    1554] = 32'hd6162f43;
    ram_cell[    1555] = 32'hcbd86d42;
    ram_cell[    1556] = 32'h577cb727;
    ram_cell[    1557] = 32'h5b843817;
    ram_cell[    1558] = 32'he3c721c3;
    ram_cell[    1559] = 32'hb2825b36;
    ram_cell[    1560] = 32'hf5e977c7;
    ram_cell[    1561] = 32'h4816f1c1;
    ram_cell[    1562] = 32'h8d6cad4e;
    ram_cell[    1563] = 32'hd57a5aee;
    ram_cell[    1564] = 32'hd70c15a9;
    ram_cell[    1565] = 32'hb6e7eaa6;
    ram_cell[    1566] = 32'h0289987d;
    ram_cell[    1567] = 32'h8e8226d0;
    ram_cell[    1568] = 32'hec05c7e0;
    ram_cell[    1569] = 32'h370c74e8;
    ram_cell[    1570] = 32'hb19be469;
    ram_cell[    1571] = 32'h7e950b96;
    ram_cell[    1572] = 32'hcb9ce546;
    ram_cell[    1573] = 32'hd529b6a3;
    ram_cell[    1574] = 32'h79a6cc64;
    ram_cell[    1575] = 32'h9eaa391f;
    ram_cell[    1576] = 32'h6e97fce4;
    ram_cell[    1577] = 32'h526da2d6;
    ram_cell[    1578] = 32'h383895a1;
    ram_cell[    1579] = 32'h981db2aa;
    ram_cell[    1580] = 32'h28b3ccb0;
    ram_cell[    1581] = 32'h09aa6dd4;
    ram_cell[    1582] = 32'h6ca24f04;
    ram_cell[    1583] = 32'hb4c620bd;
    ram_cell[    1584] = 32'h7a21678a;
    ram_cell[    1585] = 32'hcf25db67;
    ram_cell[    1586] = 32'hed7d2856;
    ram_cell[    1587] = 32'h3e311643;
    ram_cell[    1588] = 32'had802af9;
    ram_cell[    1589] = 32'h027c0dbe;
    ram_cell[    1590] = 32'h659cd6a0;
    ram_cell[    1591] = 32'hc20aa5d0;
    ram_cell[    1592] = 32'h02a1336a;
    ram_cell[    1593] = 32'hd74ce0a5;
    ram_cell[    1594] = 32'h16540ffd;
    ram_cell[    1595] = 32'h5712ffea;
    ram_cell[    1596] = 32'hf6e8e6f4;
    ram_cell[    1597] = 32'h8c4b5eb2;
    ram_cell[    1598] = 32'h2ec761de;
    ram_cell[    1599] = 32'h66d0c262;
    ram_cell[    1600] = 32'hb7b228bd;
    ram_cell[    1601] = 32'hf2860ae5;
    ram_cell[    1602] = 32'h3a9b9cee;
    ram_cell[    1603] = 32'haaa61fb2;
    ram_cell[    1604] = 32'h580c0f2c;
    ram_cell[    1605] = 32'h49b2fecf;
    ram_cell[    1606] = 32'hb96c824a;
    ram_cell[    1607] = 32'h048ff02e;
    ram_cell[    1608] = 32'h58f5d187;
    ram_cell[    1609] = 32'h28b47c3f;
    ram_cell[    1610] = 32'hd5332f5f;
    ram_cell[    1611] = 32'h79281d5c;
    ram_cell[    1612] = 32'ha91c22c4;
    ram_cell[    1613] = 32'h39f17824;
    ram_cell[    1614] = 32'h73a2c504;
    ram_cell[    1615] = 32'h22d0b8c9;
    ram_cell[    1616] = 32'hdb880ee6;
    ram_cell[    1617] = 32'ha4394616;
    ram_cell[    1618] = 32'h642e4bbc;
    ram_cell[    1619] = 32'hab767fee;
    ram_cell[    1620] = 32'haf33c9b8;
    ram_cell[    1621] = 32'h2770f7c4;
    ram_cell[    1622] = 32'hac3bef23;
    ram_cell[    1623] = 32'hd955aa19;
    ram_cell[    1624] = 32'hdafddee1;
    ram_cell[    1625] = 32'hb4d4b8c5;
    ram_cell[    1626] = 32'h9c262aed;
    ram_cell[    1627] = 32'h475d5d39;
    ram_cell[    1628] = 32'hb16b6c58;
    ram_cell[    1629] = 32'hd7b97ded;
    ram_cell[    1630] = 32'he16a5566;
    ram_cell[    1631] = 32'h8ebee3ae;
    ram_cell[    1632] = 32'h4049c366;
    ram_cell[    1633] = 32'he5bfef08;
    ram_cell[    1634] = 32'he223f0f7;
    ram_cell[    1635] = 32'h198d860a;
    ram_cell[    1636] = 32'h5572b5b5;
    ram_cell[    1637] = 32'h83ceac1c;
    ram_cell[    1638] = 32'h0a1f221f;
    ram_cell[    1639] = 32'h775b0a5f;
    ram_cell[    1640] = 32'hf4aa54f9;
    ram_cell[    1641] = 32'h565c9dd4;
    ram_cell[    1642] = 32'h490333d9;
    ram_cell[    1643] = 32'hd3790694;
    ram_cell[    1644] = 32'h88a3ac59;
    ram_cell[    1645] = 32'h389fc91e;
    ram_cell[    1646] = 32'h3c622323;
    ram_cell[    1647] = 32'h0938bbc8;
    ram_cell[    1648] = 32'hda625742;
    ram_cell[    1649] = 32'h836e5f93;
    ram_cell[    1650] = 32'h8ad21e7d;
    ram_cell[    1651] = 32'hcf1f32cd;
    ram_cell[    1652] = 32'h586591e7;
    ram_cell[    1653] = 32'h65f49a23;
    ram_cell[    1654] = 32'hd897d83f;
    ram_cell[    1655] = 32'hf7df0377;
    ram_cell[    1656] = 32'hd8a4a927;
    ram_cell[    1657] = 32'hb6438fa4;
    ram_cell[    1658] = 32'hcf075d50;
    ram_cell[    1659] = 32'hdbdbc40a;
    ram_cell[    1660] = 32'ha31ef61a;
    ram_cell[    1661] = 32'h4a322a3a;
    ram_cell[    1662] = 32'hbd04270c;
    ram_cell[    1663] = 32'h1473c66d;
    ram_cell[    1664] = 32'ha98dc4dc;
    ram_cell[    1665] = 32'hf07df272;
    ram_cell[    1666] = 32'h61ccd11e;
    ram_cell[    1667] = 32'h14b5b13d;
    ram_cell[    1668] = 32'h1a71ab47;
    ram_cell[    1669] = 32'he849bb35;
    ram_cell[    1670] = 32'h149acb59;
    ram_cell[    1671] = 32'hb3a08c29;
    ram_cell[    1672] = 32'h6c4d4a87;
    ram_cell[    1673] = 32'h2908b2f4;
    ram_cell[    1674] = 32'h684ff085;
    ram_cell[    1675] = 32'h7d4b75c5;
    ram_cell[    1676] = 32'hf04ae016;
    ram_cell[    1677] = 32'h6f910afc;
    ram_cell[    1678] = 32'ha2980618;
    ram_cell[    1679] = 32'hcf295999;
    ram_cell[    1680] = 32'h48762a50;
    ram_cell[    1681] = 32'ha96db3b1;
    ram_cell[    1682] = 32'h61bcd968;
    ram_cell[    1683] = 32'h3176767b;
    ram_cell[    1684] = 32'h9a7416f6;
    ram_cell[    1685] = 32'hf6813289;
    ram_cell[    1686] = 32'hfe08519e;
    ram_cell[    1687] = 32'h8d16d7a0;
    ram_cell[    1688] = 32'hfed0cf2a;
    ram_cell[    1689] = 32'h65f5f68d;
    ram_cell[    1690] = 32'h3ff7d801;
    ram_cell[    1691] = 32'h27610e9c;
    ram_cell[    1692] = 32'he87b0410;
    ram_cell[    1693] = 32'h3e7f7f1d;
    ram_cell[    1694] = 32'hdb1d16f5;
    ram_cell[    1695] = 32'hf7931a6b;
    ram_cell[    1696] = 32'h80c2aecc;
    ram_cell[    1697] = 32'hcf6ee0a1;
    ram_cell[    1698] = 32'ha3fa92db;
    ram_cell[    1699] = 32'hf07fcf44;
    ram_cell[    1700] = 32'h34c854ea;
    ram_cell[    1701] = 32'hce631134;
    ram_cell[    1702] = 32'hbfde4a1b;
    ram_cell[    1703] = 32'hf9e35425;
    ram_cell[    1704] = 32'hfbfc56e9;
    ram_cell[    1705] = 32'he2b4ba69;
    ram_cell[    1706] = 32'hb6b7d99a;
    ram_cell[    1707] = 32'hc6190dad;
    ram_cell[    1708] = 32'hb90d31ca;
    ram_cell[    1709] = 32'h766a861f;
    ram_cell[    1710] = 32'hdf9a572e;
    ram_cell[    1711] = 32'h33d7cbb1;
    ram_cell[    1712] = 32'hce0bd9d1;
    ram_cell[    1713] = 32'h595bb709;
    ram_cell[    1714] = 32'hde5e1176;
    ram_cell[    1715] = 32'ha69ad670;
    ram_cell[    1716] = 32'hdc3496f6;
    ram_cell[    1717] = 32'hc997cfd7;
    ram_cell[    1718] = 32'h66ccd4c0;
    ram_cell[    1719] = 32'h01001d27;
    ram_cell[    1720] = 32'ha99244e3;
    ram_cell[    1721] = 32'h4ab967d5;
    ram_cell[    1722] = 32'h597cc920;
    ram_cell[    1723] = 32'h4f52171e;
    ram_cell[    1724] = 32'h3e525dd4;
    ram_cell[    1725] = 32'hbe57bb5f;
    ram_cell[    1726] = 32'h80540ed9;
    ram_cell[    1727] = 32'h2ae919d9;
    ram_cell[    1728] = 32'h6f925323;
    ram_cell[    1729] = 32'hc49f9fa8;
    ram_cell[    1730] = 32'he9f4d067;
    ram_cell[    1731] = 32'he3fffd5d;
    ram_cell[    1732] = 32'h5e1ca1db;
    ram_cell[    1733] = 32'h4b25007f;
    ram_cell[    1734] = 32'h09263591;
    ram_cell[    1735] = 32'hfeeb6780;
    ram_cell[    1736] = 32'h287542a5;
    ram_cell[    1737] = 32'hd2b4e861;
    ram_cell[    1738] = 32'h7bf5441a;
    ram_cell[    1739] = 32'h9b4f35e7;
    ram_cell[    1740] = 32'h87c06306;
    ram_cell[    1741] = 32'h1a984ba3;
    ram_cell[    1742] = 32'h070f9251;
    ram_cell[    1743] = 32'hb69f239d;
    ram_cell[    1744] = 32'h5990fd1d;
    ram_cell[    1745] = 32'h8bf9e2b0;
    ram_cell[    1746] = 32'hcb0c055c;
    ram_cell[    1747] = 32'h40438aaf;
    ram_cell[    1748] = 32'h878abe3a;
    ram_cell[    1749] = 32'h97056995;
    ram_cell[    1750] = 32'h36d870a5;
    ram_cell[    1751] = 32'h9cd700ec;
    ram_cell[    1752] = 32'hb66eddf4;
    ram_cell[    1753] = 32'ha5d69b31;
    ram_cell[    1754] = 32'hf8891239;
    ram_cell[    1755] = 32'h7465703e;
    ram_cell[    1756] = 32'hfffb5857;
    ram_cell[    1757] = 32'h999f96ff;
    ram_cell[    1758] = 32'h16f94762;
    ram_cell[    1759] = 32'hff876018;
    ram_cell[    1760] = 32'h02e80e9f;
    ram_cell[    1761] = 32'hd67a139f;
    ram_cell[    1762] = 32'h68106393;
    ram_cell[    1763] = 32'hb8645301;
    ram_cell[    1764] = 32'hf5a93aae;
    ram_cell[    1765] = 32'h048363ab;
    ram_cell[    1766] = 32'h0518b2f3;
    ram_cell[    1767] = 32'h2726b365;
    ram_cell[    1768] = 32'hb71f141e;
    ram_cell[    1769] = 32'hdf645826;
    ram_cell[    1770] = 32'h2b37880c;
    ram_cell[    1771] = 32'h72befcec;
    ram_cell[    1772] = 32'h38585503;
    ram_cell[    1773] = 32'h467a9b4f;
    ram_cell[    1774] = 32'h47feb891;
    ram_cell[    1775] = 32'hb0d8480d;
    ram_cell[    1776] = 32'hd4caa94d;
    ram_cell[    1777] = 32'ha6171715;
    ram_cell[    1778] = 32'ha80d0d88;
    ram_cell[    1779] = 32'h99b851a7;
    ram_cell[    1780] = 32'hddbd6f21;
    ram_cell[    1781] = 32'hb91c02ef;
    ram_cell[    1782] = 32'h86691043;
    ram_cell[    1783] = 32'hcbefd027;
    ram_cell[    1784] = 32'h42e7c42b;
    ram_cell[    1785] = 32'h51e8d350;
    ram_cell[    1786] = 32'h1c136e62;
    ram_cell[    1787] = 32'ha9ee5b03;
    ram_cell[    1788] = 32'hea4b62c5;
    ram_cell[    1789] = 32'h5a5eb9f8;
    ram_cell[    1790] = 32'hd952ee8b;
    ram_cell[    1791] = 32'hcf496d59;
    ram_cell[    1792] = 32'h88b5a3eb;
    ram_cell[    1793] = 32'hd778d89a;
    ram_cell[    1794] = 32'h4a544e6f;
    ram_cell[    1795] = 32'he04a5524;
    ram_cell[    1796] = 32'hd854e372;
    ram_cell[    1797] = 32'h566cccc5;
    ram_cell[    1798] = 32'hde9f315e;
    ram_cell[    1799] = 32'h6567d108;
    ram_cell[    1800] = 32'h4160cddc;
    ram_cell[    1801] = 32'h0aeeb70e;
    ram_cell[    1802] = 32'h77daa1a7;
    ram_cell[    1803] = 32'h403a2ac9;
    ram_cell[    1804] = 32'hc75384aa;
    ram_cell[    1805] = 32'hda51aedd;
    ram_cell[    1806] = 32'hb289e239;
    ram_cell[    1807] = 32'hffc3f1f4;
    ram_cell[    1808] = 32'hc363de8f;
    ram_cell[    1809] = 32'h3d29b2bb;
    ram_cell[    1810] = 32'h4997ec7a;
    ram_cell[    1811] = 32'h5c767ad2;
    ram_cell[    1812] = 32'h4c5e63c1;
    ram_cell[    1813] = 32'h2252f6b0;
    ram_cell[    1814] = 32'h938b73c1;
    ram_cell[    1815] = 32'hb2112399;
    ram_cell[    1816] = 32'hb4d337f5;
    ram_cell[    1817] = 32'habf29359;
    ram_cell[    1818] = 32'hfe91428d;
    ram_cell[    1819] = 32'h8a9220d5;
    ram_cell[    1820] = 32'h77e08cd3;
    ram_cell[    1821] = 32'heebe4591;
    ram_cell[    1822] = 32'h44f3f8fd;
    ram_cell[    1823] = 32'h1f985929;
    ram_cell[    1824] = 32'h98c22e44;
    ram_cell[    1825] = 32'hea82cdbb;
    ram_cell[    1826] = 32'h88da9036;
    ram_cell[    1827] = 32'h6776d236;
    ram_cell[    1828] = 32'h64581170;
    ram_cell[    1829] = 32'ha487cfec;
    ram_cell[    1830] = 32'hcf4e9750;
    ram_cell[    1831] = 32'h7c4be28a;
    ram_cell[    1832] = 32'h185f8e94;
    ram_cell[    1833] = 32'hbc368776;
    ram_cell[    1834] = 32'h187735d2;
    ram_cell[    1835] = 32'h829cf162;
    ram_cell[    1836] = 32'h8c0f41ff;
    ram_cell[    1837] = 32'h3b30e715;
    ram_cell[    1838] = 32'hf609c342;
    ram_cell[    1839] = 32'hdbf70a6d;
    ram_cell[    1840] = 32'h20d4546a;
    ram_cell[    1841] = 32'h46885ff1;
    ram_cell[    1842] = 32'h456a1358;
    ram_cell[    1843] = 32'hbfb2d800;
    ram_cell[    1844] = 32'hce9bbad9;
    ram_cell[    1845] = 32'hadf00816;
    ram_cell[    1846] = 32'h235ed1fd;
    ram_cell[    1847] = 32'h3b8de44c;
    ram_cell[    1848] = 32'h24d9bfc4;
    ram_cell[    1849] = 32'h38cf2b07;
    ram_cell[    1850] = 32'h1b6ab48d;
    ram_cell[    1851] = 32'h6a8618d3;
    ram_cell[    1852] = 32'hcef49412;
    ram_cell[    1853] = 32'hb7483ca3;
    ram_cell[    1854] = 32'h2e1d033b;
    ram_cell[    1855] = 32'hdd6c6a8f;
    ram_cell[    1856] = 32'h414bb887;
    ram_cell[    1857] = 32'h06da4f9e;
    ram_cell[    1858] = 32'hf262b0fb;
    ram_cell[    1859] = 32'h95ffa053;
    ram_cell[    1860] = 32'hdd85e65a;
    ram_cell[    1861] = 32'h74c8b065;
    ram_cell[    1862] = 32'haf5820f4;
    ram_cell[    1863] = 32'h855bf15a;
    ram_cell[    1864] = 32'hf00ce716;
    ram_cell[    1865] = 32'h10322138;
    ram_cell[    1866] = 32'hf9191e65;
    ram_cell[    1867] = 32'ha23fb768;
    ram_cell[    1868] = 32'ha6a373b7;
    ram_cell[    1869] = 32'h25375070;
    ram_cell[    1870] = 32'h0191f600;
    ram_cell[    1871] = 32'h0af90504;
    ram_cell[    1872] = 32'h5a180359;
    ram_cell[    1873] = 32'hac9ec5de;
    ram_cell[    1874] = 32'h4f141b69;
    ram_cell[    1875] = 32'h986dec79;
    ram_cell[    1876] = 32'h6f2d3031;
    ram_cell[    1877] = 32'hef0bd1bf;
    ram_cell[    1878] = 32'h3075066d;
    ram_cell[    1879] = 32'hdaba9577;
    ram_cell[    1880] = 32'h2131158a;
    ram_cell[    1881] = 32'h6fdc4551;
    ram_cell[    1882] = 32'hfc3018fd;
    ram_cell[    1883] = 32'h45c4bf20;
    ram_cell[    1884] = 32'hcba2acd3;
    ram_cell[    1885] = 32'ha2176edf;
    ram_cell[    1886] = 32'h89a50233;
    ram_cell[    1887] = 32'h7e3be482;
    ram_cell[    1888] = 32'h52105f57;
    ram_cell[    1889] = 32'h1b70e26a;
    ram_cell[    1890] = 32'h2fc736bd;
    ram_cell[    1891] = 32'h59551cc0;
    ram_cell[    1892] = 32'hef56e1f0;
    ram_cell[    1893] = 32'h7b451f2c;
    ram_cell[    1894] = 32'hfe9d01a4;
    ram_cell[    1895] = 32'hcce90997;
    ram_cell[    1896] = 32'h848f6609;
    ram_cell[    1897] = 32'h973dab84;
    ram_cell[    1898] = 32'h3a59b844;
    ram_cell[    1899] = 32'ha4a77597;
    ram_cell[    1900] = 32'h11625742;
    ram_cell[    1901] = 32'hd66b523d;
    ram_cell[    1902] = 32'he41df70c;
    ram_cell[    1903] = 32'ha5c7184d;
    ram_cell[    1904] = 32'he62411fc;
    ram_cell[    1905] = 32'h142cb1f5;
    ram_cell[    1906] = 32'hc9b3180c;
    ram_cell[    1907] = 32'h59de7b68;
    ram_cell[    1908] = 32'h451abf4c;
    ram_cell[    1909] = 32'hb6e12965;
    ram_cell[    1910] = 32'h662fb481;
    ram_cell[    1911] = 32'hc150426b;
    ram_cell[    1912] = 32'h077c5b0c;
    ram_cell[    1913] = 32'hec7562aa;
    ram_cell[    1914] = 32'h8513509f;
    ram_cell[    1915] = 32'h835c37a7;
    ram_cell[    1916] = 32'h237721fb;
    ram_cell[    1917] = 32'hdeea0d0f;
    ram_cell[    1918] = 32'hffd91064;
    ram_cell[    1919] = 32'h33668110;
    ram_cell[    1920] = 32'haa76a8fb;
    ram_cell[    1921] = 32'h5bce9613;
    ram_cell[    1922] = 32'h796207d5;
    ram_cell[    1923] = 32'hc119a0b0;
    ram_cell[    1924] = 32'ha15b5886;
    ram_cell[    1925] = 32'ha7c1b012;
    ram_cell[    1926] = 32'h6c73955b;
    ram_cell[    1927] = 32'hb7824f5d;
    ram_cell[    1928] = 32'h4999f09b;
    ram_cell[    1929] = 32'h760b5f0d;
    ram_cell[    1930] = 32'h7bdfefdd;
    ram_cell[    1931] = 32'hd339f4dd;
    ram_cell[    1932] = 32'hd177ff55;
    ram_cell[    1933] = 32'he5932367;
    ram_cell[    1934] = 32'hc09b08fd;
    ram_cell[    1935] = 32'h296986c8;
    ram_cell[    1936] = 32'h3dd67c85;
    ram_cell[    1937] = 32'h7005b900;
    ram_cell[    1938] = 32'h02231589;
    ram_cell[    1939] = 32'h03d0fd5e;
    ram_cell[    1940] = 32'h6d7ac610;
    ram_cell[    1941] = 32'h6e7453a0;
    ram_cell[    1942] = 32'hf6e7c0c9;
    ram_cell[    1943] = 32'hbf3098c5;
    ram_cell[    1944] = 32'h3ef39915;
    ram_cell[    1945] = 32'hc788bffe;
    ram_cell[    1946] = 32'h329dfd40;
    ram_cell[    1947] = 32'hc4d0d52f;
    ram_cell[    1948] = 32'hdcd055f6;
    ram_cell[    1949] = 32'ha9b1ae23;
    ram_cell[    1950] = 32'hd1c59761;
    ram_cell[    1951] = 32'hde459818;
    ram_cell[    1952] = 32'hcc59d0bd;
    ram_cell[    1953] = 32'hae84d86a;
    ram_cell[    1954] = 32'h12a0929a;
    ram_cell[    1955] = 32'h7cfa6d39;
    ram_cell[    1956] = 32'h9cf9bcfa;
    ram_cell[    1957] = 32'h59e24d0d;
    ram_cell[    1958] = 32'h802a99eb;
    ram_cell[    1959] = 32'h6c336abe;
    ram_cell[    1960] = 32'h15cbbdcb;
    ram_cell[    1961] = 32'h44b6270b;
    ram_cell[    1962] = 32'h41d1b136;
    ram_cell[    1963] = 32'hdb9c64ba;
    ram_cell[    1964] = 32'h6607659f;
    ram_cell[    1965] = 32'h66a6e179;
    ram_cell[    1966] = 32'h410dc42b;
    ram_cell[    1967] = 32'hb78a0678;
    ram_cell[    1968] = 32'hc8480f5c;
    ram_cell[    1969] = 32'hfd90ea4d;
    ram_cell[    1970] = 32'h37dbc3ba;
    ram_cell[    1971] = 32'hf1814036;
    ram_cell[    1972] = 32'hfd1bbca8;
    ram_cell[    1973] = 32'h661b3a1a;
    ram_cell[    1974] = 32'h8f4d1a98;
    ram_cell[    1975] = 32'h4e600e9f;
    ram_cell[    1976] = 32'hb5a40696;
    ram_cell[    1977] = 32'h11298dda;
    ram_cell[    1978] = 32'h049f5104;
    ram_cell[    1979] = 32'he8e88ca0;
    ram_cell[    1980] = 32'h0170236e;
    ram_cell[    1981] = 32'hbe77c22d;
    ram_cell[    1982] = 32'h93d51b2c;
    ram_cell[    1983] = 32'h1fc4eb4d;
    ram_cell[    1984] = 32'h0c700ca4;
    ram_cell[    1985] = 32'hb8d0351c;
    ram_cell[    1986] = 32'h11086200;
    ram_cell[    1987] = 32'hb9675bf5;
    ram_cell[    1988] = 32'h822a3b9d;
    ram_cell[    1989] = 32'h1957ab53;
    ram_cell[    1990] = 32'hf079dedb;
    ram_cell[    1991] = 32'hee95ad3b;
    ram_cell[    1992] = 32'hd86b9e8f;
    ram_cell[    1993] = 32'h5be008fb;
    ram_cell[    1994] = 32'h90d64980;
    ram_cell[    1995] = 32'h7b638fd0;
    ram_cell[    1996] = 32'hbd424280;
    ram_cell[    1997] = 32'h3b473dac;
    ram_cell[    1998] = 32'h65d7e6c2;
    ram_cell[    1999] = 32'ha9893283;
    ram_cell[    2000] = 32'hc14923cd;
    ram_cell[    2001] = 32'h7d2176b8;
    ram_cell[    2002] = 32'ha63b9898;
    ram_cell[    2003] = 32'hd253639a;
    ram_cell[    2004] = 32'h8913d150;
    ram_cell[    2005] = 32'h4a425942;
    ram_cell[    2006] = 32'hedadb48b;
    ram_cell[    2007] = 32'h7f539465;
    ram_cell[    2008] = 32'h6f37c7cc;
    ram_cell[    2009] = 32'h4213cfab;
    ram_cell[    2010] = 32'h5b9a64e5;
    ram_cell[    2011] = 32'h3cf03072;
    ram_cell[    2012] = 32'he483efbe;
    ram_cell[    2013] = 32'h99984a4c;
    ram_cell[    2014] = 32'h13da14eb;
    ram_cell[    2015] = 32'h54adf659;
    ram_cell[    2016] = 32'ha3af9d99;
    ram_cell[    2017] = 32'hd37b1949;
    ram_cell[    2018] = 32'hf0158d02;
    ram_cell[    2019] = 32'hc6d65210;
    ram_cell[    2020] = 32'h95935107;
    ram_cell[    2021] = 32'h796f63cc;
    ram_cell[    2022] = 32'h636d5253;
    ram_cell[    2023] = 32'haed79615;
    ram_cell[    2024] = 32'ha6537981;
    ram_cell[    2025] = 32'hb3a9465c;
    ram_cell[    2026] = 32'h84ffc6d1;
    ram_cell[    2027] = 32'h052ab16c;
    ram_cell[    2028] = 32'h0ad1f898;
    ram_cell[    2029] = 32'hd96897b3;
    ram_cell[    2030] = 32'h76f97a99;
    ram_cell[    2031] = 32'hb5c20b34;
    ram_cell[    2032] = 32'h5994e682;
    ram_cell[    2033] = 32'h672ea5db;
    ram_cell[    2034] = 32'ha93d4948;
    ram_cell[    2035] = 32'h84bd64ce;
    ram_cell[    2036] = 32'h627a1ecd;
    ram_cell[    2037] = 32'hdc5e5890;
    ram_cell[    2038] = 32'h1dae73dc;
    ram_cell[    2039] = 32'hadbe8acc;
    ram_cell[    2040] = 32'h93a8182b;
    ram_cell[    2041] = 32'he0e381e2;
    ram_cell[    2042] = 32'h40cb016f;
    ram_cell[    2043] = 32'h9ba2bcc1;
    ram_cell[    2044] = 32'h26368247;
    ram_cell[    2045] = 32'h80ef25ec;
    ram_cell[    2046] = 32'h101f27b2;
    ram_cell[    2047] = 32'hb4550fc1;
    // src matrix B
    ram_cell[    2048] = 32'h106137e6;
    ram_cell[    2049] = 32'hf48d03c9;
    ram_cell[    2050] = 32'h72af95af;
    ram_cell[    2051] = 32'h324df0b2;
    ram_cell[    2052] = 32'he9728f3b;
    ram_cell[    2053] = 32'hd8214237;
    ram_cell[    2054] = 32'h329d01fe;
    ram_cell[    2055] = 32'h9fe51808;
    ram_cell[    2056] = 32'hdac96376;
    ram_cell[    2057] = 32'h4074f2df;
    ram_cell[    2058] = 32'he2126bcb;
    ram_cell[    2059] = 32'hd72140a0;
    ram_cell[    2060] = 32'h55e2d86b;
    ram_cell[    2061] = 32'h3f2043e4;
    ram_cell[    2062] = 32'h911bfe84;
    ram_cell[    2063] = 32'h8ea69ba9;
    ram_cell[    2064] = 32'h9a9f2363;
    ram_cell[    2065] = 32'ha73a01db;
    ram_cell[    2066] = 32'h866bf45a;
    ram_cell[    2067] = 32'h3df8aa4e;
    ram_cell[    2068] = 32'h5e2baff9;
    ram_cell[    2069] = 32'hfd2971c0;
    ram_cell[    2070] = 32'h2bba73aa;
    ram_cell[    2071] = 32'h99fa3fea;
    ram_cell[    2072] = 32'h599f2693;
    ram_cell[    2073] = 32'h0ad9eadc;
    ram_cell[    2074] = 32'hc84d2706;
    ram_cell[    2075] = 32'h97ecf1d4;
    ram_cell[    2076] = 32'h7a47046d;
    ram_cell[    2077] = 32'h3cbb2439;
    ram_cell[    2078] = 32'h8f82c61d;
    ram_cell[    2079] = 32'h44554e13;
    ram_cell[    2080] = 32'h23e922ed;
    ram_cell[    2081] = 32'hb5e71ba2;
    ram_cell[    2082] = 32'h9c90508b;
    ram_cell[    2083] = 32'h5c6e027d;
    ram_cell[    2084] = 32'hc060317d;
    ram_cell[    2085] = 32'hc5b3ee57;
    ram_cell[    2086] = 32'h4a72c78c;
    ram_cell[    2087] = 32'he3e64d80;
    ram_cell[    2088] = 32'hfcda6f27;
    ram_cell[    2089] = 32'h5a91bcc9;
    ram_cell[    2090] = 32'hdf04c90f;
    ram_cell[    2091] = 32'h8222b47e;
    ram_cell[    2092] = 32'h3417c5de;
    ram_cell[    2093] = 32'h51a309ac;
    ram_cell[    2094] = 32'h40e71546;
    ram_cell[    2095] = 32'h12af6cac;
    ram_cell[    2096] = 32'h44540960;
    ram_cell[    2097] = 32'h4a097e28;
    ram_cell[    2098] = 32'h1a67e29e;
    ram_cell[    2099] = 32'h0d32526b;
    ram_cell[    2100] = 32'hc58807cc;
    ram_cell[    2101] = 32'h6cf7bb7e;
    ram_cell[    2102] = 32'h454db451;
    ram_cell[    2103] = 32'hb358f801;
    ram_cell[    2104] = 32'hfcf742bc;
    ram_cell[    2105] = 32'h0c56b7f6;
    ram_cell[    2106] = 32'h7322c8dc;
    ram_cell[    2107] = 32'h04f625d6;
    ram_cell[    2108] = 32'h3872d286;
    ram_cell[    2109] = 32'h06573e04;
    ram_cell[    2110] = 32'h6ba2fc60;
    ram_cell[    2111] = 32'hff427840;
    ram_cell[    2112] = 32'heebfdc68;
    ram_cell[    2113] = 32'h29f5b6b2;
    ram_cell[    2114] = 32'h4d25607a;
    ram_cell[    2115] = 32'h20f95d53;
    ram_cell[    2116] = 32'h433795c3;
    ram_cell[    2117] = 32'h1ef4d2bf;
    ram_cell[    2118] = 32'h2fbae748;
    ram_cell[    2119] = 32'h25dce80d;
    ram_cell[    2120] = 32'h646b7f6f;
    ram_cell[    2121] = 32'hd9b98c51;
    ram_cell[    2122] = 32'h1c7b74ee;
    ram_cell[    2123] = 32'h22232b1b;
    ram_cell[    2124] = 32'h9a732f56;
    ram_cell[    2125] = 32'h4bcb277a;
    ram_cell[    2126] = 32'h7040df98;
    ram_cell[    2127] = 32'h91eab54f;
    ram_cell[    2128] = 32'h31901fcb;
    ram_cell[    2129] = 32'h3e75fbee;
    ram_cell[    2130] = 32'h270d2c14;
    ram_cell[    2131] = 32'hd9fb84b7;
    ram_cell[    2132] = 32'h327218e2;
    ram_cell[    2133] = 32'h08631586;
    ram_cell[    2134] = 32'hc81df348;
    ram_cell[    2135] = 32'h1e51a777;
    ram_cell[    2136] = 32'h0d38fbfb;
    ram_cell[    2137] = 32'h9fd0d37c;
    ram_cell[    2138] = 32'h71255b07;
    ram_cell[    2139] = 32'h51ae9e73;
    ram_cell[    2140] = 32'he10b9304;
    ram_cell[    2141] = 32'h0836613d;
    ram_cell[    2142] = 32'h1d0624f9;
    ram_cell[    2143] = 32'h6217594d;
    ram_cell[    2144] = 32'h23294d4d;
    ram_cell[    2145] = 32'hca01c322;
    ram_cell[    2146] = 32'heb3daa63;
    ram_cell[    2147] = 32'h5b008ae3;
    ram_cell[    2148] = 32'h45e3ca67;
    ram_cell[    2149] = 32'h8f46c6a8;
    ram_cell[    2150] = 32'h0573c625;
    ram_cell[    2151] = 32'h1f5b1b00;
    ram_cell[    2152] = 32'hbc19667b;
    ram_cell[    2153] = 32'ha45d41d0;
    ram_cell[    2154] = 32'h6769702f;
    ram_cell[    2155] = 32'h62272e63;
    ram_cell[    2156] = 32'hae91c17c;
    ram_cell[    2157] = 32'h9a03b269;
    ram_cell[    2158] = 32'h21ad2b65;
    ram_cell[    2159] = 32'h8faa6515;
    ram_cell[    2160] = 32'h9d423173;
    ram_cell[    2161] = 32'h6a50d8f6;
    ram_cell[    2162] = 32'h2a103cf0;
    ram_cell[    2163] = 32'h4da8a622;
    ram_cell[    2164] = 32'h1c5c77bc;
    ram_cell[    2165] = 32'h08ed1617;
    ram_cell[    2166] = 32'hcec010e9;
    ram_cell[    2167] = 32'h8c1324c4;
    ram_cell[    2168] = 32'h7cddca91;
    ram_cell[    2169] = 32'h12043cab;
    ram_cell[    2170] = 32'h1a9c5587;
    ram_cell[    2171] = 32'ha9bd89e5;
    ram_cell[    2172] = 32'h4f980ee0;
    ram_cell[    2173] = 32'h8a914adb;
    ram_cell[    2174] = 32'hf5a83ef2;
    ram_cell[    2175] = 32'h82621f79;
    ram_cell[    2176] = 32'h8f26ffad;
    ram_cell[    2177] = 32'hc55b1445;
    ram_cell[    2178] = 32'h6f8998a9;
    ram_cell[    2179] = 32'h69b42cea;
    ram_cell[    2180] = 32'haf114e25;
    ram_cell[    2181] = 32'hb1605e96;
    ram_cell[    2182] = 32'h65d7e1a3;
    ram_cell[    2183] = 32'hba2a9db8;
    ram_cell[    2184] = 32'h20bcf6f5;
    ram_cell[    2185] = 32'hb372d3c9;
    ram_cell[    2186] = 32'hc0848f00;
    ram_cell[    2187] = 32'h1ae9cf40;
    ram_cell[    2188] = 32'h14058f7f;
    ram_cell[    2189] = 32'hb150c69c;
    ram_cell[    2190] = 32'hf88b2618;
    ram_cell[    2191] = 32'h23ef5dd5;
    ram_cell[    2192] = 32'h12c8d108;
    ram_cell[    2193] = 32'hff7b0c47;
    ram_cell[    2194] = 32'h2786e82a;
    ram_cell[    2195] = 32'h3d616b69;
    ram_cell[    2196] = 32'h7efdaa6b;
    ram_cell[    2197] = 32'h75a13279;
    ram_cell[    2198] = 32'h20a58d32;
    ram_cell[    2199] = 32'h5dde405f;
    ram_cell[    2200] = 32'hd1455960;
    ram_cell[    2201] = 32'h63cdc325;
    ram_cell[    2202] = 32'h56cce3c1;
    ram_cell[    2203] = 32'h628670b6;
    ram_cell[    2204] = 32'he3cf6885;
    ram_cell[    2205] = 32'h7c4771bc;
    ram_cell[    2206] = 32'hcedb6808;
    ram_cell[    2207] = 32'hdb7a9c22;
    ram_cell[    2208] = 32'hc26eaa1d;
    ram_cell[    2209] = 32'h9e2cae5e;
    ram_cell[    2210] = 32'hb131b766;
    ram_cell[    2211] = 32'h7d135128;
    ram_cell[    2212] = 32'h020b962e;
    ram_cell[    2213] = 32'h539ad4d6;
    ram_cell[    2214] = 32'he2ee1e3b;
    ram_cell[    2215] = 32'hb8e1462a;
    ram_cell[    2216] = 32'h6830dcd3;
    ram_cell[    2217] = 32'h735ff7a9;
    ram_cell[    2218] = 32'hf7e04c48;
    ram_cell[    2219] = 32'hccac1537;
    ram_cell[    2220] = 32'h9e1a920f;
    ram_cell[    2221] = 32'hecc1a1ce;
    ram_cell[    2222] = 32'h72ce453d;
    ram_cell[    2223] = 32'h9fd46ee9;
    ram_cell[    2224] = 32'h3ccd7f3c;
    ram_cell[    2225] = 32'h639742ee;
    ram_cell[    2226] = 32'h03a30fe9;
    ram_cell[    2227] = 32'h15522161;
    ram_cell[    2228] = 32'ha21c50fb;
    ram_cell[    2229] = 32'h45445b56;
    ram_cell[    2230] = 32'h1bbb0246;
    ram_cell[    2231] = 32'h2083e078;
    ram_cell[    2232] = 32'hb9d2827b;
    ram_cell[    2233] = 32'hf322ced1;
    ram_cell[    2234] = 32'hb0604458;
    ram_cell[    2235] = 32'h73e74b33;
    ram_cell[    2236] = 32'h5befd2e1;
    ram_cell[    2237] = 32'h14cf3109;
    ram_cell[    2238] = 32'h82316ed9;
    ram_cell[    2239] = 32'hc9355adc;
    ram_cell[    2240] = 32'h93a05374;
    ram_cell[    2241] = 32'h87b2d31b;
    ram_cell[    2242] = 32'had7e19ff;
    ram_cell[    2243] = 32'h0b119493;
    ram_cell[    2244] = 32'h1f6c890c;
    ram_cell[    2245] = 32'h11019324;
    ram_cell[    2246] = 32'hc119c23e;
    ram_cell[    2247] = 32'h549a9f1f;
    ram_cell[    2248] = 32'h2994680b;
    ram_cell[    2249] = 32'h1d54079d;
    ram_cell[    2250] = 32'h712488d9;
    ram_cell[    2251] = 32'h8f06d7db;
    ram_cell[    2252] = 32'h980e9fa5;
    ram_cell[    2253] = 32'ha9ddea65;
    ram_cell[    2254] = 32'h2eef5902;
    ram_cell[    2255] = 32'h4990e796;
    ram_cell[    2256] = 32'hff437c01;
    ram_cell[    2257] = 32'h8124bdb8;
    ram_cell[    2258] = 32'hb24c1ce7;
    ram_cell[    2259] = 32'h1e797501;
    ram_cell[    2260] = 32'hdbd5c520;
    ram_cell[    2261] = 32'hf8349283;
    ram_cell[    2262] = 32'hf7af2e5c;
    ram_cell[    2263] = 32'h6ec4cc0b;
    ram_cell[    2264] = 32'he0be6139;
    ram_cell[    2265] = 32'h951be53b;
    ram_cell[    2266] = 32'hf604d769;
    ram_cell[    2267] = 32'hebca9b7f;
    ram_cell[    2268] = 32'h0d3aad39;
    ram_cell[    2269] = 32'h286048ea;
    ram_cell[    2270] = 32'hd0f669e7;
    ram_cell[    2271] = 32'h13e867b2;
    ram_cell[    2272] = 32'h28226186;
    ram_cell[    2273] = 32'hc4452679;
    ram_cell[    2274] = 32'h7c2d69c4;
    ram_cell[    2275] = 32'h90bddb44;
    ram_cell[    2276] = 32'hf22797c8;
    ram_cell[    2277] = 32'hd5a99cb5;
    ram_cell[    2278] = 32'hf124ac52;
    ram_cell[    2279] = 32'h792d7f3f;
    ram_cell[    2280] = 32'h1a95d27d;
    ram_cell[    2281] = 32'h85d7ea34;
    ram_cell[    2282] = 32'h28135aef;
    ram_cell[    2283] = 32'h1fc85402;
    ram_cell[    2284] = 32'h625ecaca;
    ram_cell[    2285] = 32'h34c51a6e;
    ram_cell[    2286] = 32'hbeba6bfa;
    ram_cell[    2287] = 32'h4caad662;
    ram_cell[    2288] = 32'h9b60f655;
    ram_cell[    2289] = 32'h276727ac;
    ram_cell[    2290] = 32'h28a450e6;
    ram_cell[    2291] = 32'h86a42c6a;
    ram_cell[    2292] = 32'h44ffc723;
    ram_cell[    2293] = 32'h83e8df47;
    ram_cell[    2294] = 32'h0e9b96d6;
    ram_cell[    2295] = 32'h67d36825;
    ram_cell[    2296] = 32'h5795d98d;
    ram_cell[    2297] = 32'h72524d85;
    ram_cell[    2298] = 32'h44072c6a;
    ram_cell[    2299] = 32'he9ef5806;
    ram_cell[    2300] = 32'hc260ce11;
    ram_cell[    2301] = 32'hfd82ba4f;
    ram_cell[    2302] = 32'ha3cda24a;
    ram_cell[    2303] = 32'h6a542e89;
    ram_cell[    2304] = 32'h2ecd7285;
    ram_cell[    2305] = 32'hb60c0d9d;
    ram_cell[    2306] = 32'h93d26820;
    ram_cell[    2307] = 32'h67f1b696;
    ram_cell[    2308] = 32'h798e36e0;
    ram_cell[    2309] = 32'he9be9f88;
    ram_cell[    2310] = 32'ha8460570;
    ram_cell[    2311] = 32'h968d82cc;
    ram_cell[    2312] = 32'hf4c422b4;
    ram_cell[    2313] = 32'h2b4209e2;
    ram_cell[    2314] = 32'h1a3e2350;
    ram_cell[    2315] = 32'hdfdf058f;
    ram_cell[    2316] = 32'h5b785d6c;
    ram_cell[    2317] = 32'h2a6b93f0;
    ram_cell[    2318] = 32'ha3c5aca4;
    ram_cell[    2319] = 32'he9740879;
    ram_cell[    2320] = 32'hccf1ad24;
    ram_cell[    2321] = 32'h775a71d8;
    ram_cell[    2322] = 32'hc9035cdb;
    ram_cell[    2323] = 32'hab00990f;
    ram_cell[    2324] = 32'h0b987f2b;
    ram_cell[    2325] = 32'h04d0756c;
    ram_cell[    2326] = 32'h067ea87c;
    ram_cell[    2327] = 32'h21499611;
    ram_cell[    2328] = 32'h3196db67;
    ram_cell[    2329] = 32'h3449e9f3;
    ram_cell[    2330] = 32'h952e74fe;
    ram_cell[    2331] = 32'h63c7bd73;
    ram_cell[    2332] = 32'h201d2cd5;
    ram_cell[    2333] = 32'he419c0fa;
    ram_cell[    2334] = 32'h097c4d55;
    ram_cell[    2335] = 32'hbd7d59b2;
    ram_cell[    2336] = 32'h39edcf06;
    ram_cell[    2337] = 32'h97dd149e;
    ram_cell[    2338] = 32'h938b010f;
    ram_cell[    2339] = 32'h06867a21;
    ram_cell[    2340] = 32'h7eed501b;
    ram_cell[    2341] = 32'h92b00eb3;
    ram_cell[    2342] = 32'h7f97f7e1;
    ram_cell[    2343] = 32'hd7418534;
    ram_cell[    2344] = 32'h56abd247;
    ram_cell[    2345] = 32'h1ac87865;
    ram_cell[    2346] = 32'h77189cc4;
    ram_cell[    2347] = 32'h8a4ca67f;
    ram_cell[    2348] = 32'h3044d0d3;
    ram_cell[    2349] = 32'h5465cf15;
    ram_cell[    2350] = 32'h8dc070d7;
    ram_cell[    2351] = 32'h279ec4b7;
    ram_cell[    2352] = 32'h2afa009b;
    ram_cell[    2353] = 32'h8e604b56;
    ram_cell[    2354] = 32'h154143a8;
    ram_cell[    2355] = 32'h1b1b0aeb;
    ram_cell[    2356] = 32'he5eb25a8;
    ram_cell[    2357] = 32'h991a0b02;
    ram_cell[    2358] = 32'hf2fdadca;
    ram_cell[    2359] = 32'hc946e5fe;
    ram_cell[    2360] = 32'hfce58b7c;
    ram_cell[    2361] = 32'h9eeadb3a;
    ram_cell[    2362] = 32'h73744fd3;
    ram_cell[    2363] = 32'h08669e46;
    ram_cell[    2364] = 32'h08851bd4;
    ram_cell[    2365] = 32'h238b2ded;
    ram_cell[    2366] = 32'h86308248;
    ram_cell[    2367] = 32'hdd20d31e;
    ram_cell[    2368] = 32'h174ab19b;
    ram_cell[    2369] = 32'h6a9d2345;
    ram_cell[    2370] = 32'h505f6892;
    ram_cell[    2371] = 32'h9970caa7;
    ram_cell[    2372] = 32'h5be579b8;
    ram_cell[    2373] = 32'h57f92949;
    ram_cell[    2374] = 32'h1a22c67c;
    ram_cell[    2375] = 32'h8c2b7427;
    ram_cell[    2376] = 32'h46d73c2a;
    ram_cell[    2377] = 32'h139f25c3;
    ram_cell[    2378] = 32'h3c60cf86;
    ram_cell[    2379] = 32'haab9afcb;
    ram_cell[    2380] = 32'h8e6779b5;
    ram_cell[    2381] = 32'h0fc14e4a;
    ram_cell[    2382] = 32'hb202063c;
    ram_cell[    2383] = 32'h713b23e0;
    ram_cell[    2384] = 32'h65b882a8;
    ram_cell[    2385] = 32'ha4014812;
    ram_cell[    2386] = 32'h7ad719a1;
    ram_cell[    2387] = 32'h293d34a4;
    ram_cell[    2388] = 32'hb89a38dc;
    ram_cell[    2389] = 32'hd222bab8;
    ram_cell[    2390] = 32'h86687ded;
    ram_cell[    2391] = 32'h40fa8cea;
    ram_cell[    2392] = 32'h26cdf350;
    ram_cell[    2393] = 32'h2f008aae;
    ram_cell[    2394] = 32'h7841588f;
    ram_cell[    2395] = 32'hf781ffc0;
    ram_cell[    2396] = 32'h16c029e2;
    ram_cell[    2397] = 32'hc97304e6;
    ram_cell[    2398] = 32'h1874333a;
    ram_cell[    2399] = 32'hf2cf46f5;
    ram_cell[    2400] = 32'h1964f92d;
    ram_cell[    2401] = 32'hb94fe465;
    ram_cell[    2402] = 32'h2776f0d4;
    ram_cell[    2403] = 32'hf66bf03f;
    ram_cell[    2404] = 32'h568b9e65;
    ram_cell[    2405] = 32'h927512de;
    ram_cell[    2406] = 32'ha4f63a8a;
    ram_cell[    2407] = 32'h9657fca5;
    ram_cell[    2408] = 32'h7e4a5d93;
    ram_cell[    2409] = 32'h9e483932;
    ram_cell[    2410] = 32'ha280daa0;
    ram_cell[    2411] = 32'h91e2e4f6;
    ram_cell[    2412] = 32'h83f8ae5f;
    ram_cell[    2413] = 32'h0aec5cb3;
    ram_cell[    2414] = 32'hd3564f3a;
    ram_cell[    2415] = 32'hcbd9da42;
    ram_cell[    2416] = 32'hd906f097;
    ram_cell[    2417] = 32'h5d0ecc60;
    ram_cell[    2418] = 32'h513ab73d;
    ram_cell[    2419] = 32'h76b3cf80;
    ram_cell[    2420] = 32'h0254f2a3;
    ram_cell[    2421] = 32'h82934038;
    ram_cell[    2422] = 32'h09d3ae44;
    ram_cell[    2423] = 32'hf37b56e4;
    ram_cell[    2424] = 32'hc3b633dd;
    ram_cell[    2425] = 32'ha5f3e682;
    ram_cell[    2426] = 32'hacd15cc5;
    ram_cell[    2427] = 32'h83307a72;
    ram_cell[    2428] = 32'h7a69515c;
    ram_cell[    2429] = 32'h68b27933;
    ram_cell[    2430] = 32'hb8973d0b;
    ram_cell[    2431] = 32'hce3289c1;
    ram_cell[    2432] = 32'ha5098585;
    ram_cell[    2433] = 32'hcf4a28dd;
    ram_cell[    2434] = 32'h1b34a633;
    ram_cell[    2435] = 32'h18cd31d9;
    ram_cell[    2436] = 32'h6f7e75f3;
    ram_cell[    2437] = 32'h8af02e48;
    ram_cell[    2438] = 32'hb0963f4c;
    ram_cell[    2439] = 32'h36042d20;
    ram_cell[    2440] = 32'h8d086138;
    ram_cell[    2441] = 32'he1f50b83;
    ram_cell[    2442] = 32'h28406a7f;
    ram_cell[    2443] = 32'h03182d55;
    ram_cell[    2444] = 32'h3a4e0e44;
    ram_cell[    2445] = 32'h9565b4fc;
    ram_cell[    2446] = 32'h27d12d6e;
    ram_cell[    2447] = 32'hc14f8b3f;
    ram_cell[    2448] = 32'h95efbe0e;
    ram_cell[    2449] = 32'h79a676a1;
    ram_cell[    2450] = 32'hb4726241;
    ram_cell[    2451] = 32'hc2f91c01;
    ram_cell[    2452] = 32'h917cd3de;
    ram_cell[    2453] = 32'h6af76dd0;
    ram_cell[    2454] = 32'he51252e1;
    ram_cell[    2455] = 32'h82c04254;
    ram_cell[    2456] = 32'he17def0e;
    ram_cell[    2457] = 32'h4018fbca;
    ram_cell[    2458] = 32'hae30bbb8;
    ram_cell[    2459] = 32'h3b0fd325;
    ram_cell[    2460] = 32'h4576cf87;
    ram_cell[    2461] = 32'h99ce6537;
    ram_cell[    2462] = 32'h89d6f3ae;
    ram_cell[    2463] = 32'h3b9a4aa1;
    ram_cell[    2464] = 32'h31da089c;
    ram_cell[    2465] = 32'h88454788;
    ram_cell[    2466] = 32'h20124fdc;
    ram_cell[    2467] = 32'hf446e856;
    ram_cell[    2468] = 32'hbc064a1a;
    ram_cell[    2469] = 32'h3f4eb091;
    ram_cell[    2470] = 32'hae080741;
    ram_cell[    2471] = 32'hd6984437;
    ram_cell[    2472] = 32'he08a9e34;
    ram_cell[    2473] = 32'h3f91a7a4;
    ram_cell[    2474] = 32'h5fd2eb00;
    ram_cell[    2475] = 32'h081ef2ca;
    ram_cell[    2476] = 32'hd9312f00;
    ram_cell[    2477] = 32'h3f00f756;
    ram_cell[    2478] = 32'hc70bbf5a;
    ram_cell[    2479] = 32'he39f898a;
    ram_cell[    2480] = 32'heaf03033;
    ram_cell[    2481] = 32'had4ff47d;
    ram_cell[    2482] = 32'h75ffe469;
    ram_cell[    2483] = 32'h008b69d1;
    ram_cell[    2484] = 32'hcc1afd3e;
    ram_cell[    2485] = 32'h83d022c6;
    ram_cell[    2486] = 32'h189c5a50;
    ram_cell[    2487] = 32'h54dc6ff6;
    ram_cell[    2488] = 32'h6f616560;
    ram_cell[    2489] = 32'h72d7b0a4;
    ram_cell[    2490] = 32'hd1a222d8;
    ram_cell[    2491] = 32'h06ec91d5;
    ram_cell[    2492] = 32'h509cf3e6;
    ram_cell[    2493] = 32'h711fe58d;
    ram_cell[    2494] = 32'hce0d26d2;
    ram_cell[    2495] = 32'h15feed9d;
    ram_cell[    2496] = 32'h1a6d7440;
    ram_cell[    2497] = 32'h1a9306a2;
    ram_cell[    2498] = 32'h52a81f40;
    ram_cell[    2499] = 32'h72a0a7e8;
    ram_cell[    2500] = 32'h7a780120;
    ram_cell[    2501] = 32'hcb3360ca;
    ram_cell[    2502] = 32'he20dcbbb;
    ram_cell[    2503] = 32'h1c785966;
    ram_cell[    2504] = 32'h09249dd5;
    ram_cell[    2505] = 32'h2a448814;
    ram_cell[    2506] = 32'hbf9ab218;
    ram_cell[    2507] = 32'h99b93886;
    ram_cell[    2508] = 32'h02c6ddb7;
    ram_cell[    2509] = 32'h342facee;
    ram_cell[    2510] = 32'hf0121c38;
    ram_cell[    2511] = 32'h4165eeb7;
    ram_cell[    2512] = 32'h386d2586;
    ram_cell[    2513] = 32'h0bb51a0b;
    ram_cell[    2514] = 32'h7ef7ca1c;
    ram_cell[    2515] = 32'he077c1a8;
    ram_cell[    2516] = 32'h4b0f2475;
    ram_cell[    2517] = 32'hbe123f9e;
    ram_cell[    2518] = 32'h2c12d34f;
    ram_cell[    2519] = 32'h4d3d90ed;
    ram_cell[    2520] = 32'h2d7d1d37;
    ram_cell[    2521] = 32'he3f95f11;
    ram_cell[    2522] = 32'h7d274df4;
    ram_cell[    2523] = 32'hc609d8a0;
    ram_cell[    2524] = 32'hdd23d63a;
    ram_cell[    2525] = 32'h48e9a7de;
    ram_cell[    2526] = 32'h55b124b3;
    ram_cell[    2527] = 32'h529aba2d;
    ram_cell[    2528] = 32'h1d1bf870;
    ram_cell[    2529] = 32'h7fcd0068;
    ram_cell[    2530] = 32'h663b1ee3;
    ram_cell[    2531] = 32'h64aff900;
    ram_cell[    2532] = 32'h8a9737eb;
    ram_cell[    2533] = 32'hedd802aa;
    ram_cell[    2534] = 32'h27c24ca6;
    ram_cell[    2535] = 32'h6dfddbb8;
    ram_cell[    2536] = 32'h3ce25d12;
    ram_cell[    2537] = 32'h83c22931;
    ram_cell[    2538] = 32'hd10d4fc9;
    ram_cell[    2539] = 32'h421fb27f;
    ram_cell[    2540] = 32'h1bcf0686;
    ram_cell[    2541] = 32'h80abaeba;
    ram_cell[    2542] = 32'hbcc7d2b4;
    ram_cell[    2543] = 32'hc3cfe0a0;
    ram_cell[    2544] = 32'h69401510;
    ram_cell[    2545] = 32'h70d85369;
    ram_cell[    2546] = 32'h9fed477c;
    ram_cell[    2547] = 32'hee310627;
    ram_cell[    2548] = 32'hc7046245;
    ram_cell[    2549] = 32'h81378de7;
    ram_cell[    2550] = 32'ha2b177ba;
    ram_cell[    2551] = 32'hf5d5a45a;
    ram_cell[    2552] = 32'h17f4fc76;
    ram_cell[    2553] = 32'hf02a3321;
    ram_cell[    2554] = 32'h62b4b1fc;
    ram_cell[    2555] = 32'h0421147a;
    ram_cell[    2556] = 32'he7376e3f;
    ram_cell[    2557] = 32'hd5888eb9;
    ram_cell[    2558] = 32'h09efc225;
    ram_cell[    2559] = 32'h93355adf;
    ram_cell[    2560] = 32'h05349c46;
    ram_cell[    2561] = 32'h0c7b3528;
    ram_cell[    2562] = 32'h815d6f5e;
    ram_cell[    2563] = 32'h2068f5c8;
    ram_cell[    2564] = 32'h7a53886c;
    ram_cell[    2565] = 32'haaa7a120;
    ram_cell[    2566] = 32'hb67f3015;
    ram_cell[    2567] = 32'hc13ffd64;
    ram_cell[    2568] = 32'h591766ec;
    ram_cell[    2569] = 32'h3b9d5980;
    ram_cell[    2570] = 32'h289279cc;
    ram_cell[    2571] = 32'hd509c7e8;
    ram_cell[    2572] = 32'hd1c528c3;
    ram_cell[    2573] = 32'hf6a9f7bd;
    ram_cell[    2574] = 32'h8bfd4413;
    ram_cell[    2575] = 32'hb238f4fc;
    ram_cell[    2576] = 32'h72acf088;
    ram_cell[    2577] = 32'hc657a4f9;
    ram_cell[    2578] = 32'hd00a2747;
    ram_cell[    2579] = 32'h7532838f;
    ram_cell[    2580] = 32'h9b6db0a6;
    ram_cell[    2581] = 32'hae7e2e54;
    ram_cell[    2582] = 32'hfef624cd;
    ram_cell[    2583] = 32'hfdaf51a7;
    ram_cell[    2584] = 32'h5a0cfcf5;
    ram_cell[    2585] = 32'h3ba0c67c;
    ram_cell[    2586] = 32'hf78e83c9;
    ram_cell[    2587] = 32'hd3f94ed4;
    ram_cell[    2588] = 32'h403652a3;
    ram_cell[    2589] = 32'h8c83618f;
    ram_cell[    2590] = 32'hcf25f7a8;
    ram_cell[    2591] = 32'h570b2f04;
    ram_cell[    2592] = 32'hb759f8f8;
    ram_cell[    2593] = 32'h86b7d38e;
    ram_cell[    2594] = 32'h96474a56;
    ram_cell[    2595] = 32'hd71f0927;
    ram_cell[    2596] = 32'h298d2613;
    ram_cell[    2597] = 32'h9722f9bf;
    ram_cell[    2598] = 32'h504ea936;
    ram_cell[    2599] = 32'h30b6a63d;
    ram_cell[    2600] = 32'hec688179;
    ram_cell[    2601] = 32'h53a3c7e0;
    ram_cell[    2602] = 32'h59438466;
    ram_cell[    2603] = 32'h1057dadb;
    ram_cell[    2604] = 32'hd6a3b121;
    ram_cell[    2605] = 32'he718e642;
    ram_cell[    2606] = 32'he9dbcc64;
    ram_cell[    2607] = 32'h2d670d3a;
    ram_cell[    2608] = 32'hfc240d90;
    ram_cell[    2609] = 32'hefe214c8;
    ram_cell[    2610] = 32'h4855e3e8;
    ram_cell[    2611] = 32'hdd3ccf81;
    ram_cell[    2612] = 32'h291f6a6e;
    ram_cell[    2613] = 32'h56422a40;
    ram_cell[    2614] = 32'h73e97076;
    ram_cell[    2615] = 32'h11b8f3fb;
    ram_cell[    2616] = 32'h49342cd6;
    ram_cell[    2617] = 32'h2b692563;
    ram_cell[    2618] = 32'h6a64d86d;
    ram_cell[    2619] = 32'h17f9ad5c;
    ram_cell[    2620] = 32'h0af5b7ae;
    ram_cell[    2621] = 32'h44e3f97b;
    ram_cell[    2622] = 32'h92b5adba;
    ram_cell[    2623] = 32'hdbc0f465;
    ram_cell[    2624] = 32'h5d297ce0;
    ram_cell[    2625] = 32'ha2ef935b;
    ram_cell[    2626] = 32'h1b953214;
    ram_cell[    2627] = 32'h1870180d;
    ram_cell[    2628] = 32'h3fb7a837;
    ram_cell[    2629] = 32'h453bd077;
    ram_cell[    2630] = 32'hbb2d0c6d;
    ram_cell[    2631] = 32'hf87dfc4c;
    ram_cell[    2632] = 32'h6496cc8a;
    ram_cell[    2633] = 32'h4b0ffd01;
    ram_cell[    2634] = 32'had6415b4;
    ram_cell[    2635] = 32'hc3e4c6c4;
    ram_cell[    2636] = 32'he91804c8;
    ram_cell[    2637] = 32'hc8080b8c;
    ram_cell[    2638] = 32'h6ec88171;
    ram_cell[    2639] = 32'hebc0841c;
    ram_cell[    2640] = 32'h4c0587b0;
    ram_cell[    2641] = 32'h905ad8ea;
    ram_cell[    2642] = 32'h1bbbc7b9;
    ram_cell[    2643] = 32'h79f5e2b6;
    ram_cell[    2644] = 32'h23e039b9;
    ram_cell[    2645] = 32'h97e575a3;
    ram_cell[    2646] = 32'hd2930aac;
    ram_cell[    2647] = 32'h0ae77922;
    ram_cell[    2648] = 32'h37105ab5;
    ram_cell[    2649] = 32'hacaac2c0;
    ram_cell[    2650] = 32'h223274ba;
    ram_cell[    2651] = 32'h2076da40;
    ram_cell[    2652] = 32'he10c7614;
    ram_cell[    2653] = 32'h19a9d55b;
    ram_cell[    2654] = 32'he605d50a;
    ram_cell[    2655] = 32'h5dfcb5c0;
    ram_cell[    2656] = 32'ha48f1c20;
    ram_cell[    2657] = 32'h92eae4ea;
    ram_cell[    2658] = 32'hd97600cd;
    ram_cell[    2659] = 32'haa54a8f7;
    ram_cell[    2660] = 32'hc22f20d4;
    ram_cell[    2661] = 32'h57778886;
    ram_cell[    2662] = 32'h2ded1bd2;
    ram_cell[    2663] = 32'h7b8d1e4f;
    ram_cell[    2664] = 32'hf8726dea;
    ram_cell[    2665] = 32'h4d84d0c6;
    ram_cell[    2666] = 32'h618348ab;
    ram_cell[    2667] = 32'h87001516;
    ram_cell[    2668] = 32'hf745c1db;
    ram_cell[    2669] = 32'h72490d3c;
    ram_cell[    2670] = 32'he0189162;
    ram_cell[    2671] = 32'h6b2338ec;
    ram_cell[    2672] = 32'h76ef8f9c;
    ram_cell[    2673] = 32'hfbd530c0;
    ram_cell[    2674] = 32'ha219c5d5;
    ram_cell[    2675] = 32'hd68d6eef;
    ram_cell[    2676] = 32'h428c3d03;
    ram_cell[    2677] = 32'h39db894b;
    ram_cell[    2678] = 32'h3d0eb343;
    ram_cell[    2679] = 32'h4610d489;
    ram_cell[    2680] = 32'h95625163;
    ram_cell[    2681] = 32'h714d668c;
    ram_cell[    2682] = 32'h3b534457;
    ram_cell[    2683] = 32'hd93b8c8c;
    ram_cell[    2684] = 32'h5006b538;
    ram_cell[    2685] = 32'h638a7621;
    ram_cell[    2686] = 32'hb153284a;
    ram_cell[    2687] = 32'h7e5f0ab1;
    ram_cell[    2688] = 32'h0f50bec7;
    ram_cell[    2689] = 32'h44daf632;
    ram_cell[    2690] = 32'h7f235c03;
    ram_cell[    2691] = 32'h5fb436ac;
    ram_cell[    2692] = 32'hc094c4eb;
    ram_cell[    2693] = 32'h101bb8d7;
    ram_cell[    2694] = 32'h2b459a08;
    ram_cell[    2695] = 32'h76e40897;
    ram_cell[    2696] = 32'hc876c989;
    ram_cell[    2697] = 32'h90594b94;
    ram_cell[    2698] = 32'hfa5b1b75;
    ram_cell[    2699] = 32'h01f62145;
    ram_cell[    2700] = 32'h82246657;
    ram_cell[    2701] = 32'hb3777317;
    ram_cell[    2702] = 32'h54282238;
    ram_cell[    2703] = 32'ha8ba6766;
    ram_cell[    2704] = 32'h4bf5cbda;
    ram_cell[    2705] = 32'hefad0e46;
    ram_cell[    2706] = 32'ha9ed588b;
    ram_cell[    2707] = 32'he2e16576;
    ram_cell[    2708] = 32'ha3147f64;
    ram_cell[    2709] = 32'h06a6e72f;
    ram_cell[    2710] = 32'h7d48410b;
    ram_cell[    2711] = 32'h1d8a40d6;
    ram_cell[    2712] = 32'hf756ab3c;
    ram_cell[    2713] = 32'h712bcc2c;
    ram_cell[    2714] = 32'hbebde368;
    ram_cell[    2715] = 32'hb0bc8510;
    ram_cell[    2716] = 32'h70639f3a;
    ram_cell[    2717] = 32'hcf87cb14;
    ram_cell[    2718] = 32'h483d8170;
    ram_cell[    2719] = 32'h5c90bf56;
    ram_cell[    2720] = 32'h0a206d4a;
    ram_cell[    2721] = 32'h8b8a5b20;
    ram_cell[    2722] = 32'h90378210;
    ram_cell[    2723] = 32'ha9854bcb;
    ram_cell[    2724] = 32'h20379a9b;
    ram_cell[    2725] = 32'hff65aadd;
    ram_cell[    2726] = 32'h3c74f22f;
    ram_cell[    2727] = 32'h7d96f2e7;
    ram_cell[    2728] = 32'h1549898e;
    ram_cell[    2729] = 32'h0c9567f7;
    ram_cell[    2730] = 32'hf60fbfbd;
    ram_cell[    2731] = 32'h68b3590e;
    ram_cell[    2732] = 32'h962d38f7;
    ram_cell[    2733] = 32'h45c2f32c;
    ram_cell[    2734] = 32'hf2febc3b;
    ram_cell[    2735] = 32'hf4a319f1;
    ram_cell[    2736] = 32'hc21d653e;
    ram_cell[    2737] = 32'h554ae000;
    ram_cell[    2738] = 32'h3ed868b9;
    ram_cell[    2739] = 32'h19dc0353;
    ram_cell[    2740] = 32'h6b3f32af;
    ram_cell[    2741] = 32'hb441e8d0;
    ram_cell[    2742] = 32'hbc9cdd2c;
    ram_cell[    2743] = 32'h9e9671a1;
    ram_cell[    2744] = 32'h2fa6b862;
    ram_cell[    2745] = 32'h1eec10dc;
    ram_cell[    2746] = 32'h81dc4cc7;
    ram_cell[    2747] = 32'h703c265c;
    ram_cell[    2748] = 32'hef875f3e;
    ram_cell[    2749] = 32'hfd6ea874;
    ram_cell[    2750] = 32'ha8f8431b;
    ram_cell[    2751] = 32'he56d5e26;
    ram_cell[    2752] = 32'h95032118;
    ram_cell[    2753] = 32'h8483b983;
    ram_cell[    2754] = 32'he80440e6;
    ram_cell[    2755] = 32'h28b19624;
    ram_cell[    2756] = 32'hd59dd1db;
    ram_cell[    2757] = 32'hf9585111;
    ram_cell[    2758] = 32'h0baa1cea;
    ram_cell[    2759] = 32'h8100dc4b;
    ram_cell[    2760] = 32'h4e916dd2;
    ram_cell[    2761] = 32'hfda0f340;
    ram_cell[    2762] = 32'hd4ebcfe6;
    ram_cell[    2763] = 32'haf19ed4e;
    ram_cell[    2764] = 32'h56725c37;
    ram_cell[    2765] = 32'he8331044;
    ram_cell[    2766] = 32'h8f287230;
    ram_cell[    2767] = 32'h03c442ec;
    ram_cell[    2768] = 32'h0fe28450;
    ram_cell[    2769] = 32'hfc63c999;
    ram_cell[    2770] = 32'h2d5a3e24;
    ram_cell[    2771] = 32'h61467db7;
    ram_cell[    2772] = 32'h67b7b747;
    ram_cell[    2773] = 32'head3588f;
    ram_cell[    2774] = 32'h9887e746;
    ram_cell[    2775] = 32'hc7822549;
    ram_cell[    2776] = 32'hf22bbbfb;
    ram_cell[    2777] = 32'hbae44367;
    ram_cell[    2778] = 32'hfc546ead;
    ram_cell[    2779] = 32'h8725d22f;
    ram_cell[    2780] = 32'had4c2edb;
    ram_cell[    2781] = 32'h449d5da7;
    ram_cell[    2782] = 32'hf906092b;
    ram_cell[    2783] = 32'h69d1bc3e;
    ram_cell[    2784] = 32'h3d8d5746;
    ram_cell[    2785] = 32'h1898f504;
    ram_cell[    2786] = 32'h49adbdb1;
    ram_cell[    2787] = 32'haac5600b;
    ram_cell[    2788] = 32'hc982bef2;
    ram_cell[    2789] = 32'h3f23fb1e;
    ram_cell[    2790] = 32'ha445d7f3;
    ram_cell[    2791] = 32'hc2724c7d;
    ram_cell[    2792] = 32'hd2b25cd4;
    ram_cell[    2793] = 32'h839da74b;
    ram_cell[    2794] = 32'h5141555f;
    ram_cell[    2795] = 32'ha79116f7;
    ram_cell[    2796] = 32'h86800406;
    ram_cell[    2797] = 32'hd9bfd3d6;
    ram_cell[    2798] = 32'he3f356e1;
    ram_cell[    2799] = 32'h892213cf;
    ram_cell[    2800] = 32'hcf47dda7;
    ram_cell[    2801] = 32'h02946697;
    ram_cell[    2802] = 32'h6a79260e;
    ram_cell[    2803] = 32'hc450351c;
    ram_cell[    2804] = 32'hd374d16d;
    ram_cell[    2805] = 32'h7229a185;
    ram_cell[    2806] = 32'hbeee1717;
    ram_cell[    2807] = 32'hc197c639;
    ram_cell[    2808] = 32'h5462b4a4;
    ram_cell[    2809] = 32'hcd9149d7;
    ram_cell[    2810] = 32'h041d571f;
    ram_cell[    2811] = 32'ha4c02b9e;
    ram_cell[    2812] = 32'h9dc9cb53;
    ram_cell[    2813] = 32'h640a6f43;
    ram_cell[    2814] = 32'hb9715811;
    ram_cell[    2815] = 32'hf22fe463;
    ram_cell[    2816] = 32'h211996b0;
    ram_cell[    2817] = 32'hd82246ae;
    ram_cell[    2818] = 32'h4e1d7291;
    ram_cell[    2819] = 32'hedd97aea;
    ram_cell[    2820] = 32'h09f0c32b;
    ram_cell[    2821] = 32'h76f722ad;
    ram_cell[    2822] = 32'h65c58121;
    ram_cell[    2823] = 32'h363bdac7;
    ram_cell[    2824] = 32'h3792062e;
    ram_cell[    2825] = 32'h6556021a;
    ram_cell[    2826] = 32'hbe12d0ee;
    ram_cell[    2827] = 32'hf3977344;
    ram_cell[    2828] = 32'h2b4e24c4;
    ram_cell[    2829] = 32'hccaca29e;
    ram_cell[    2830] = 32'hf3bfe1ba;
    ram_cell[    2831] = 32'h9c9bf91a;
    ram_cell[    2832] = 32'hae5e6aeb;
    ram_cell[    2833] = 32'h53c7a37c;
    ram_cell[    2834] = 32'h602a9063;
    ram_cell[    2835] = 32'h2ff66363;
    ram_cell[    2836] = 32'h14d46652;
    ram_cell[    2837] = 32'h9c658106;
    ram_cell[    2838] = 32'he81435e1;
    ram_cell[    2839] = 32'h0444cad5;
    ram_cell[    2840] = 32'hae70533d;
    ram_cell[    2841] = 32'hfddbcc55;
    ram_cell[    2842] = 32'ha1607418;
    ram_cell[    2843] = 32'h3621b977;
    ram_cell[    2844] = 32'h4600b9ad;
    ram_cell[    2845] = 32'h10a6b3ca;
    ram_cell[    2846] = 32'hbc02118a;
    ram_cell[    2847] = 32'h24bb7a00;
    ram_cell[    2848] = 32'hb30b3736;
    ram_cell[    2849] = 32'h53e1dbe5;
    ram_cell[    2850] = 32'hbaed7cc0;
    ram_cell[    2851] = 32'haed7742c;
    ram_cell[    2852] = 32'h6a79311d;
    ram_cell[    2853] = 32'h7b5cb7db;
    ram_cell[    2854] = 32'h59880a4b;
    ram_cell[    2855] = 32'h2f303606;
    ram_cell[    2856] = 32'h5797e996;
    ram_cell[    2857] = 32'hd038b00d;
    ram_cell[    2858] = 32'hb7ae9cec;
    ram_cell[    2859] = 32'hf8ec1eb2;
    ram_cell[    2860] = 32'h930ad90f;
    ram_cell[    2861] = 32'hd059eac7;
    ram_cell[    2862] = 32'hfb4f4cf3;
    ram_cell[    2863] = 32'h0adfe024;
    ram_cell[    2864] = 32'h017e2fb1;
    ram_cell[    2865] = 32'hfe67eb83;
    ram_cell[    2866] = 32'hb5e48010;
    ram_cell[    2867] = 32'h82a365aa;
    ram_cell[    2868] = 32'h66799e42;
    ram_cell[    2869] = 32'h3d57fd5f;
    ram_cell[    2870] = 32'h5419396a;
    ram_cell[    2871] = 32'h2aa3b2fe;
    ram_cell[    2872] = 32'h97c3635f;
    ram_cell[    2873] = 32'h879b5a67;
    ram_cell[    2874] = 32'hb02d6fa3;
    ram_cell[    2875] = 32'hbbd3ccd9;
    ram_cell[    2876] = 32'h28ddd3eb;
    ram_cell[    2877] = 32'hf391dce0;
    ram_cell[    2878] = 32'hb23eec64;
    ram_cell[    2879] = 32'h0f711670;
    ram_cell[    2880] = 32'h17e92482;
    ram_cell[    2881] = 32'ha45deea7;
    ram_cell[    2882] = 32'hb8431d73;
    ram_cell[    2883] = 32'h810bb270;
    ram_cell[    2884] = 32'h6e02c739;
    ram_cell[    2885] = 32'h9f919fd8;
    ram_cell[    2886] = 32'h6a51d421;
    ram_cell[    2887] = 32'h9c9fb597;
    ram_cell[    2888] = 32'h00dc8e08;
    ram_cell[    2889] = 32'hba1b59bb;
    ram_cell[    2890] = 32'he5e26d31;
    ram_cell[    2891] = 32'h90b6efa5;
    ram_cell[    2892] = 32'he59b6f3b;
    ram_cell[    2893] = 32'ha420e185;
    ram_cell[    2894] = 32'h21539255;
    ram_cell[    2895] = 32'h02a42816;
    ram_cell[    2896] = 32'ha07aa9cb;
    ram_cell[    2897] = 32'h7d991295;
    ram_cell[    2898] = 32'h811d6334;
    ram_cell[    2899] = 32'h295cd7b7;
    ram_cell[    2900] = 32'hf2d0f80f;
    ram_cell[    2901] = 32'h334de655;
    ram_cell[    2902] = 32'hd8dac81c;
    ram_cell[    2903] = 32'h7088fe66;
    ram_cell[    2904] = 32'h1a0c52ac;
    ram_cell[    2905] = 32'heebd9177;
    ram_cell[    2906] = 32'h61905bd0;
    ram_cell[    2907] = 32'hbd005342;
    ram_cell[    2908] = 32'h48374a8e;
    ram_cell[    2909] = 32'h53a9ae73;
    ram_cell[    2910] = 32'h3b81ab0a;
    ram_cell[    2911] = 32'h6b762e75;
    ram_cell[    2912] = 32'he9b4cd24;
    ram_cell[    2913] = 32'h3b44b0ae;
    ram_cell[    2914] = 32'h3b328c35;
    ram_cell[    2915] = 32'h03923e83;
    ram_cell[    2916] = 32'h4dba9937;
    ram_cell[    2917] = 32'h5c128142;
    ram_cell[    2918] = 32'h5d6677d3;
    ram_cell[    2919] = 32'h2e2ac979;
    ram_cell[    2920] = 32'h2a61fd1b;
    ram_cell[    2921] = 32'h4f272928;
    ram_cell[    2922] = 32'hddbbfe55;
    ram_cell[    2923] = 32'h68dfb8bf;
    ram_cell[    2924] = 32'ha122386c;
    ram_cell[    2925] = 32'h8fce64ec;
    ram_cell[    2926] = 32'h74e6e748;
    ram_cell[    2927] = 32'he262af67;
    ram_cell[    2928] = 32'h4f7231d3;
    ram_cell[    2929] = 32'heca2ee5f;
    ram_cell[    2930] = 32'hc12454d4;
    ram_cell[    2931] = 32'h4a66c414;
    ram_cell[    2932] = 32'hadf14b55;
    ram_cell[    2933] = 32'h65774ecc;
    ram_cell[    2934] = 32'hd4d1279c;
    ram_cell[    2935] = 32'h9db5e91a;
    ram_cell[    2936] = 32'hc6aacbc0;
    ram_cell[    2937] = 32'he355ad8f;
    ram_cell[    2938] = 32'hc7bbe340;
    ram_cell[    2939] = 32'hb0d16c63;
    ram_cell[    2940] = 32'h22d7bf6d;
    ram_cell[    2941] = 32'h2d2eab3c;
    ram_cell[    2942] = 32'h4f9c7de7;
    ram_cell[    2943] = 32'h153178d1;
    ram_cell[    2944] = 32'h903cecac;
    ram_cell[    2945] = 32'hdaf6838c;
    ram_cell[    2946] = 32'h0b967271;
    ram_cell[    2947] = 32'h86c565bc;
    ram_cell[    2948] = 32'h38cc56bf;
    ram_cell[    2949] = 32'h703b9730;
    ram_cell[    2950] = 32'h50f77feb;
    ram_cell[    2951] = 32'hdd746096;
    ram_cell[    2952] = 32'hb1987eee;
    ram_cell[    2953] = 32'h19a4d931;
    ram_cell[    2954] = 32'hce5ef629;
    ram_cell[    2955] = 32'h6ac627b7;
    ram_cell[    2956] = 32'h07d1157a;
    ram_cell[    2957] = 32'h3eeddc69;
    ram_cell[    2958] = 32'h90e0654f;
    ram_cell[    2959] = 32'h2ff94cfd;
    ram_cell[    2960] = 32'h0e050d08;
    ram_cell[    2961] = 32'ha45184d0;
    ram_cell[    2962] = 32'h39e24ea8;
    ram_cell[    2963] = 32'hbb9b5ace;
    ram_cell[    2964] = 32'hbbdeeede;
    ram_cell[    2965] = 32'h68ef5cb9;
    ram_cell[    2966] = 32'h4ffa30ce;
    ram_cell[    2967] = 32'hbf3d8349;
    ram_cell[    2968] = 32'h846bd117;
    ram_cell[    2969] = 32'h429cacff;
    ram_cell[    2970] = 32'ha5688f70;
    ram_cell[    2971] = 32'ha1074d96;
    ram_cell[    2972] = 32'h9814958f;
    ram_cell[    2973] = 32'h835b84f4;
    ram_cell[    2974] = 32'h98c000f1;
    ram_cell[    2975] = 32'h1965cd88;
    ram_cell[    2976] = 32'hf60a9e3b;
    ram_cell[    2977] = 32'h645b9c28;
    ram_cell[    2978] = 32'hf6d4c85c;
    ram_cell[    2979] = 32'hbe1ab941;
    ram_cell[    2980] = 32'hd6ab9a4b;
    ram_cell[    2981] = 32'ha0734805;
    ram_cell[    2982] = 32'hfe8d7172;
    ram_cell[    2983] = 32'hdc44604f;
    ram_cell[    2984] = 32'h354357c5;
    ram_cell[    2985] = 32'h46b457c5;
    ram_cell[    2986] = 32'h128cc052;
    ram_cell[    2987] = 32'he4b3cd75;
    ram_cell[    2988] = 32'hf7f54adf;
    ram_cell[    2989] = 32'h76ce4376;
    ram_cell[    2990] = 32'hdcf4b07d;
    ram_cell[    2991] = 32'h8c26a88b;
    ram_cell[    2992] = 32'hba97a261;
    ram_cell[    2993] = 32'h3a49c3d4;
    ram_cell[    2994] = 32'h491e4d81;
    ram_cell[    2995] = 32'h16c3f24f;
    ram_cell[    2996] = 32'he8196251;
    ram_cell[    2997] = 32'hf478266d;
    ram_cell[    2998] = 32'ha9b219b6;
    ram_cell[    2999] = 32'ha7587e66;
    ram_cell[    3000] = 32'h1285378f;
    ram_cell[    3001] = 32'h93f80c57;
    ram_cell[    3002] = 32'hefb83c8c;
    ram_cell[    3003] = 32'ha9da98f5;
    ram_cell[    3004] = 32'hfd331c70;
    ram_cell[    3005] = 32'h3d42fb1c;
    ram_cell[    3006] = 32'he2018f3d;
    ram_cell[    3007] = 32'h4d33d67c;
    ram_cell[    3008] = 32'hcfe4458c;
    ram_cell[    3009] = 32'ha43f2340;
    ram_cell[    3010] = 32'h0430ae46;
    ram_cell[    3011] = 32'h6f801f05;
    ram_cell[    3012] = 32'h6a2b3d3f;
    ram_cell[    3013] = 32'h726998cc;
    ram_cell[    3014] = 32'hed6ee2bf;
    ram_cell[    3015] = 32'h6db0bf43;
    ram_cell[    3016] = 32'hf64d5c37;
    ram_cell[    3017] = 32'hebf50268;
    ram_cell[    3018] = 32'hf6db1a4d;
    ram_cell[    3019] = 32'ha69be425;
    ram_cell[    3020] = 32'hf1ff8f00;
    ram_cell[    3021] = 32'hb29c6e2c;
    ram_cell[    3022] = 32'h2ac045df;
    ram_cell[    3023] = 32'hf239f640;
    ram_cell[    3024] = 32'h5264f46b;
    ram_cell[    3025] = 32'h1e1d2133;
    ram_cell[    3026] = 32'hd340e3d7;
    ram_cell[    3027] = 32'h93c3eb67;
    ram_cell[    3028] = 32'ha08fb593;
    ram_cell[    3029] = 32'hc4787996;
    ram_cell[    3030] = 32'hc4377ad5;
    ram_cell[    3031] = 32'h0a86d97a;
    ram_cell[    3032] = 32'hcaecacaa;
    ram_cell[    3033] = 32'h46a05832;
    ram_cell[    3034] = 32'he1e90364;
    ram_cell[    3035] = 32'h1ce2a829;
    ram_cell[    3036] = 32'h44e4fdad;
    ram_cell[    3037] = 32'h3b773f2e;
    ram_cell[    3038] = 32'hd73c1821;
    ram_cell[    3039] = 32'h7a30b341;
    ram_cell[    3040] = 32'hed853942;
    ram_cell[    3041] = 32'h3ff6a2cd;
    ram_cell[    3042] = 32'h9e441b4a;
    ram_cell[    3043] = 32'h0bad7709;
    ram_cell[    3044] = 32'h99dede61;
    ram_cell[    3045] = 32'ha8c68397;
    ram_cell[    3046] = 32'h6c9199f3;
    ram_cell[    3047] = 32'h5574cc1f;
    ram_cell[    3048] = 32'h09fccb60;
    ram_cell[    3049] = 32'ha2f36b67;
    ram_cell[    3050] = 32'hdf7f40d2;
    ram_cell[    3051] = 32'h786f7513;
    ram_cell[    3052] = 32'h7c142292;
    ram_cell[    3053] = 32'habe30b82;
    ram_cell[    3054] = 32'ha2d0d00b;
    ram_cell[    3055] = 32'hb01e6417;
    ram_cell[    3056] = 32'h9f0fea4e;
    ram_cell[    3057] = 32'h8e365d08;
    ram_cell[    3058] = 32'h26c224e4;
    ram_cell[    3059] = 32'h664086b4;
    ram_cell[    3060] = 32'ha0c77cbe;
    ram_cell[    3061] = 32'h630ad961;
    ram_cell[    3062] = 32'h9722bef6;
    ram_cell[    3063] = 32'h1b9c7322;
    ram_cell[    3064] = 32'h11f2a00c;
    ram_cell[    3065] = 32'h28dd0ae4;
    ram_cell[    3066] = 32'hb3a3cdd2;
    ram_cell[    3067] = 32'h3e11f804;
    ram_cell[    3068] = 32'hfc9389ea;
    ram_cell[    3069] = 32'h40084a54;
    ram_cell[    3070] = 32'hf833ff9e;
    ram_cell[    3071] = 32'hd427025c;
end

endmodule

